/*
 
 Conway's Game of Life modeled in SVerilog
 
 */

module datapath (clk, grid_evolve, initial_state, run, reset);

logic [255:0] 	grid;
input logic clk;
input logic [255:0]  initial_state;
input logic          reset;
input logic          run;
output logic [255:0] grid_evolve;

typedef enum 	logic [1:0] {S0, S1, S2, S3} statetype;
   statetype state, nextstate;
   
   // state register
   always_ff @(posedge clk, posedge reset)
     if (reset) state <= S0;
     else if (run) state <= S1;
     else state <= S2;
   
   // next state logic
   evolve efga (grid, grid_evolve);
   always_comb
     case (state)
       S0: begin 
         grid = initial_state;
         if(run) nextstate <= S1;
         else nextstate <= S0;
       end

       S1: begin
         grid = grid_evolve;
         if(run) nextstate <= S1;
         else if(run == 0) nextstate <= S2;
         else nextstate <= S0;
       end

       S2: begin
         if(run) nextstate <= S1;
         else if(run == 0) nextstate <= S2;
         else nextstate <= S0;
       end

       S3: begin
         nextstate <= S0;
       end
     endcase

endmodule

module evolve (grid, grid_evolve);
input logic [255:0] 	grid;
output logic [255:0] 	grid_evolve;
//row 1  
evolve3 e0 (grid_evolve[0], grid[1], grid[16], grid[17], grid[0]);
evolve5 e1 (grid_evolve[1], grid[0], grid[2], grid[16], grid[17], grid[18], grid[1]);
evolve5 e2 (grid_evolve[2], grid[1], grid[3], grid[17], grid[18], grid[19], grid[2]);
evolve5 e3 (grid_evolve[3], grid[2], grid[4], grid[18], grid[19], grid[20], grid[3]);
evolve5 e4 (grid_evolve[4], grid[3], grid[5], grid[19], grid[20], grid[21], grid[4]);
evolve5 e5 (grid_evolve[5], grid[4], grid[6], grid[20], grid[21], grid[22], grid[5]);
evolve5 e6 (grid_evolve[6], grid[5], grid[7], grid[21], grid[22], grid[23], grid[6]);
evolve5 e7 (grid_evolve[7], grid[6], grid[8], grid[22], grid[23], grid[24], grid[7]);
evolve5 e8 (grid_evolve[8], grid[7], grid[9], grid[23], grid[24], grid[25], grid[8]);
evolve5 e9 (grid_evolve[9], grid[8], grid[10], grid[24], grid[25], grid[26], grid[9]);
evolve5 e10 (grid_evolve[10], grid[9], grid[11], grid[25], grid[26], grid[27], grid[10]);
evolve5 e11 (grid_evolve[11], grid[10], grid[12], grid[26], grid[27], grid[28], grid[11]);
evolve5 e12 (grid_evolve[12], grid[11], grid[13], grid[27], grid[28], grid[29], grid[12]);
evolve5 e13 (grid_evolve[13], grid[12], grid[14], grid[28], grid[29], grid[30], grid[13]);
evolve5 e14 (grid_evolve[14], grid[13], grid[15], grid[29], grid[30], grid[31], grid[14]);
evolve3 e15 (grid_evolve[15], grid[14], grid[30], grid[31], grid[15]);

//row 2
evolve5 e16 (grid_evolve[16], grid[0], grid[1], grid[17], grid[32], grid[33], grid[16]);
evolve8 e17 (grid_evolve[17], grid[0], grid[1], grid[2], grid[16], grid[18], grid[32], grid[33], grid[34], grid[17]);
evolve8 e18 (grid_evolve[18], grid[1], grid[2], grid[3], grid[17], grid[19], grid[33], grid[34], grid[35], grid[18]);
evolve8 e19 (grid_evolve[19], grid[2], grid[3], grid[4], grid[18], grid[20], grid[34], grid[35], grid[36], grid[19]);
evolve8 e20 (grid_evolve[20], grid[3], grid[4], grid[5], grid[19], grid[21], grid[35], grid[36], grid[37], grid[20]);
evolve8 e21 (grid_evolve[21], grid[4], grid[5], grid[6], grid[20], grid[22], grid[36], grid[37], grid[38], grid[21]);
evolve8 e22 (grid_evolve[22], grid[5], grid[6], grid[7], grid[21], grid[23], grid[37], grid[38], grid[39], grid[22]);
evolve8 e23 (grid_evolve[23], grid[6], grid[7], grid[8], grid[22], grid[24], grid[38], grid[39], grid[40], grid[23]);
evolve8 e24 (grid_evolve[24], grid[7], grid[8], grid[9], grid[23], grid[25], grid[39], grid[40], grid[41], grid[24]);
evolve8 e25 (grid_evolve[25], grid[8], grid[9], grid[10], grid[24], grid[26], grid[40], grid[41], grid[42], grid[25]);
evolve8 e26 (grid_evolve[26], grid[9], grid[10], grid[11], grid[25], grid[27], grid[41], grid[42], grid[43], grid[26]);
evolve8 e27 (grid_evolve[27], grid[10], grid[11], grid[12], grid[26], grid[28], grid[42], grid[43], grid[44], grid[27]);
evolve8 e28 (grid_evolve[28], grid[11], grid[12], grid[13], grid[27], grid[29], grid[43], grid[44], grid[45], grid[28]);
evolve8 e29 (grid_evolve[29], grid[12], grid[13], grid[14], grid[28], grid[30], grid[44], grid[45], grid[46], grid[29]);
evolve8 e30 (grid_evolve[30], grid[13], grid[14], grid[15], grid[29], grid[31], grid[45], grid[46], grid[47], grid[30]);
evolve5 e31 (grid_evolve[31], grid[14], grid[15], grid[30], grid[46], grid[47], grid[31]);

//row 3
evolve5 e32 (grid_evolve[32], grid[16], grid[17], grid[33], grid[48], grid[49], grid[32]);
evolve8 e33 (grid_evolve[33], grid[16], grid[17], grid[18], grid[32], grid[34], grid[48], grid[49], grid[50], grid[33]);
evolve8 e34 (grid_evolve[34], grid[17], grid[18], grid[19], grid[33], grid[35], grid[49], grid[50], grid[51], grid[34]);
evolve8 e35 (grid_evolve[35], grid[18], grid[19], grid[20], grid[34], grid[36], grid[50], grid[51], grid[52], grid[35]);
evolve8 e36 (grid_evolve[36], grid[19], grid[20], grid[21], grid[35], grid[37], grid[51], grid[52], grid[53], grid[36]);
evolve8 e37 (grid_evolve[37], grid[20], grid[21], grid[22], grid[36], grid[38], grid[52], grid[53], grid[54], grid[37]);
evolve8 e38 (grid_evolve[38], grid[21], grid[22], grid[23], grid[37], grid[39], grid[53], grid[54], grid[55], grid[38]);
evolve8 e39 (grid_evolve[39], grid[22], grid[23], grid[24], grid[38], grid[40], grid[54], grid[55], grid[56], grid[39]);
evolve8 e40 (grid_evolve[40], grid[23], grid[24], grid[25], grid[39], grid[41], grid[55], grid[56], grid[57], grid[40]);
evolve8 e41 (grid_evolve[41], grid[24], grid[25], grid[26], grid[40], grid[42], grid[56], grid[57], grid[58], grid[41]);
evolve8 e42 (grid_evolve[42], grid[25], grid[26], grid[27], grid[41], grid[43], grid[57], grid[58], grid[59], grid[42]);
evolve8 e43 (grid_evolve[43], grid[26], grid[27], grid[28], grid[42], grid[44], grid[58], grid[59], grid[60], grid[43]);
evolve8 e44 (grid_evolve[44], grid[27], grid[28], grid[29], grid[43], grid[45], grid[59], grid[60], grid[61], grid[44]);
evolve8 e45 (grid_evolve[45], grid[28], grid[29], grid[30], grid[44], grid[46], grid[60], grid[61], grid[62], grid[45]);
evolve8 e46 (grid_evolve[46], grid[29], grid[30], grid[31], grid[45], grid[47], grid[61], grid[62], grid[63], grid[46]);
evolve5 e47 (grid_evolve[47], grid[30], grid[31], grid[46], grid[62], grid[63], grid[47]);

//row 4
evolve5 e48 (grid_evolve[48], grid[32], grid[33], grid[49], grid[64], grid[65], grid[48]);
evolve8 e49 (grid_evolve[49], grid[32], grid[33], grid[34], grid[48], grid[50], grid[64], grid[65], grid[66], grid[49]);
evolve8 e50 (grid_evolve[50], grid[33], grid[34], grid[35], grid[49], grid[51], grid[65], grid[66], grid[67], grid[50]);
evolve8 e51 (grid_evolve[51], grid[34], grid[35], grid[36], grid[50], grid[52], grid[66], grid[67], grid[68], grid[51]);
evolve8 e52 (grid_evolve[52], grid[35], grid[36], grid[37], grid[51], grid[53], grid[67], grid[68], grid[69], grid[52]);
evolve8 e53 (grid_evolve[53], grid[36], grid[37], grid[38], grid[52], grid[54], grid[68], grid[69], grid[70], grid[53]);
evolve8 e54 (grid_evolve[54], grid[37], grid[38], grid[39], grid[53], grid[55], grid[69], grid[70], grid[71], grid[54]);
evolve8 e55 (grid_evolve[55], grid[38], grid[39], grid[40], grid[54], grid[56], grid[70], grid[71], grid[72], grid[55]);
evolve8 e56 (grid_evolve[56], grid[39], grid[40], grid[41], grid[55], grid[57], grid[71], grid[72], grid[73], grid[56]);
evolve8 e57 (grid_evolve[57], grid[40], grid[41], grid[42], grid[56], grid[58], grid[72], grid[73], grid[74], grid[57]);
evolve8 e58 (grid_evolve[58], grid[41], grid[42], grid[43], grid[57], grid[59], grid[73], grid[74], grid[75], grid[58]);
evolve8 e59 (grid_evolve[59], grid[42], grid[43], grid[44], grid[58], grid[60], grid[74], grid[75], grid[76], grid[59]);
evolve8 e60 (grid_evolve[60], grid[43], grid[44], grid[45], grid[59], grid[61], grid[75], grid[76], grid[77], grid[60]);
evolve8 e61 (grid_evolve[61], grid[44], grid[45], grid[46], grid[60], grid[62], grid[76], grid[77], grid[78], grid[61]);
evolve8 e62 (grid_evolve[62], grid[45], grid[46], grid[47], grid[61], grid[63], grid[77], grid[78], grid[79], grid[62]);
evolve5 e63 (grid_evolve[63], grid[46], grid[47], grid[62], grid[78], grid[79], grid[63]);

//row 5
evolve5 e64 (grid_evolve[64], grid[48], grid[49], grid[65], grid[80], grid[81], grid[64]);
evolve8 e65 (grid_evolve[65], grid[48], grid[49], grid[50], grid[64], grid[66], grid[80], grid[81], grid[82], grid[65]);
evolve8 e66 (grid_evolve[66], grid[49], grid[50], grid[51], grid[65], grid[67], grid[81], grid[82], grid[83], grid[66]);
evolve8 e67 (grid_evolve[67], grid[50], grid[51], grid[52], grid[66], grid[68], grid[82], grid[83], grid[84], grid[67]);
evolve8 e68 (grid_evolve[68], grid[51], grid[52], grid[53], grid[67], grid[69], grid[83], grid[84], grid[85], grid[68]);
evolve8 e69 (grid_evolve[69], grid[52], grid[53], grid[54], grid[68], grid[70], grid[84], grid[85], grid[86], grid[69]);
evolve8 e70 (grid_evolve[70], grid[53], grid[54], grid[55], grid[69], grid[71], grid[85], grid[86], grid[87], grid[70]);
evolve8 e71 (grid_evolve[71], grid[54], grid[55], grid[56], grid[70], grid[72], grid[86], grid[87], grid[88], grid[71]);
evolve8 e72 (grid_evolve[72], grid[55], grid[56], grid[57], grid[71], grid[73], grid[87], grid[88], grid[89], grid[72]);
evolve8 e73 (grid_evolve[73], grid[56], grid[57], grid[58], grid[72], grid[74], grid[88], grid[89], grid[90], grid[73]);
evolve8 e74 (grid_evolve[74], grid[57], grid[58], grid[59], grid[73], grid[75], grid[89], grid[90], grid[91], grid[74]);
evolve8 e75 (grid_evolve[75], grid[58], grid[59], grid[60], grid[74], grid[76], grid[90], grid[91], grid[92], grid[75]);
evolve8 e76 (grid_evolve[76], grid[59], grid[60], grid[61], grid[75], grid[77], grid[91], grid[92], grid[93], grid[76]);
evolve8 e77 (grid_evolve[77], grid[60], grid[61], grid[62], grid[76], grid[78], grid[92], grid[93], grid[94], grid[77]);
evolve8 e78 (grid_evolve[78], grid[61], grid[62], grid[63], grid[77], grid[79], grid[93], grid[94], grid[95], grid[78]);
evolve5 e79 (grid_evolve[79], grid[62], grid[63], grid[78], grid[94], grid[95], grid[79]);

//row 6
evolve5 e80 (grid_evolve[80], grid[64], grid[65], grid[81], grid[96], grid[97], grid[80]);
evolve8 e81 (grid_evolve[81], grid[64], grid[65], grid[66], grid[80], grid[82], grid[96], grid[97], grid[98], grid[81]);
evolve8 e82 (grid_evolve[82], grid[65], grid[66], grid[67], grid[81], grid[83], grid[97], grid[98], grid[99], grid[82]);
evolve8 e83 (grid_evolve[83], grid[66], grid[67], grid[68], grid[82], grid[84], grid[98], grid[99], grid[100], grid[83]);
evolve8 e84 (grid_evolve[84], grid[67], grid[68], grid[69], grid[83], grid[85], grid[99], grid[100], grid[101], grid[84]);
evolve8 e85 (grid_evolve[85], grid[68], grid[69], grid[70], grid[84], grid[86], grid[100], grid[101], grid[102], grid[85]);
evolve8 e86 (grid_evolve[86], grid[69], grid[70], grid[71], grid[85], grid[87], grid[101], grid[102], grid[103], grid[86]);
evolve8 e87 (grid_evolve[87], grid[70], grid[71], grid[72], grid[86], grid[88], grid[102], grid[103], grid[104], grid[87]);
evolve8 e88 (grid_evolve[88], grid[71], grid[72], grid[73], grid[87], grid[89], grid[103], grid[104], grid[105], grid[88]);
evolve8 e89 (grid_evolve[89], grid[72], grid[73], grid[74], grid[88], grid[90], grid[104], grid[105], grid[106], grid[89]);
evolve8 e90 (grid_evolve[90], grid[73], grid[74], grid[75], grid[89], grid[91], grid[105], grid[106], grid[107], grid[90]);
evolve8 e91 (grid_evolve[91], grid[74], grid[75], grid[76], grid[90], grid[92], grid[106], grid[107], grid[108], grid[91]);
evolve8 e92 (grid_evolve[92], grid[75], grid[76], grid[77], grid[91], grid[93], grid[107], grid[108], grid[109], grid[92]);
evolve8 e93 (grid_evolve[93], grid[76], grid[77], grid[78], grid[92], grid[94], grid[108], grid[109], grid[110], grid[93]);
evolve8 e94 (grid_evolve[94], grid[77], grid[78], grid[79], grid[93], grid[95], grid[109], grid[110], grid[111], grid[94]);
evolve5 e95 (grid_evolve[95], grid[78], grid[79], grid[94], grid[110], grid[111], grid[95]);

//row 7
evolve5 e96 (grid_evolve[96], grid[80], grid[81], grid[97], grid[112], grid[113], grid[96]);
evolve8 e97 (grid_evolve[97], grid[80], grid[81], grid[82], grid[96], grid[98], grid[112], grid[113], grid[114], grid[97]);
evolve8 e98 (grid_evolve[98], grid[81], grid[82], grid[83], grid[97], grid[99], grid[113], grid[114], grid[115], grid[98]);
evolve8 e99 (grid_evolve[99], grid[82], grid[83], grid[84], grid[98], grid[100], grid[114], grid[115], grid[116], grid[99]);
evolve8 e100 (grid_evolve[100], grid[83], grid[84], grid[85], grid[99], grid[101], grid[115], grid[116], grid[117], grid[100]);
evolve8 e101 (grid_evolve[101], grid[84], grid[85], grid[86], grid[100], grid[102], grid[116], grid[117], grid[118], grid[101]);
evolve8 e102 (grid_evolve[102], grid[85], grid[86], grid[87], grid[101], grid[103], grid[117], grid[118], grid[119], grid[102]);
evolve8 e103 (grid_evolve[103], grid[86], grid[87], grid[88], grid[102], grid[104], grid[118], grid[119], grid[120], grid[103]);
evolve8 e104 (grid_evolve[104], grid[87], grid[88], grid[89], grid[103], grid[105], grid[119], grid[120], grid[121], grid[104]);
evolve8 e105 (grid_evolve[105], grid[88], grid[89], grid[90], grid[104], grid[106], grid[120], grid[121], grid[122], grid[105]);
evolve8 e106 (grid_evolve[106], grid[89], grid[90], grid[91], grid[105], grid[107], grid[121], grid[122], grid[123], grid[106]);
evolve8 e107 (grid_evolve[107], grid[90], grid[91], grid[92], grid[106], grid[108], grid[122], grid[123], grid[124], grid[107]);
evolve8 e108 (grid_evolve[108], grid[91], grid[92], grid[93], grid[107], grid[109], grid[123], grid[124], grid[125], grid[108]);
evolve8 e109 (grid_evolve[109], grid[92], grid[93], grid[94], grid[108], grid[110], grid[124], grid[125], grid[126], grid[109]);
evolve8 e110 (grid_evolve[110], grid[93], grid[94], grid[95], grid[109], grid[111], grid[125], grid[126], grid[127], grid[110]);
evolve5 e111 (grid_evolve[111], grid[94], grid[95], grid[110], grid[126], grid[127], grid[111]);

//row 8
evolve5 e112 (grid_evolve[112], grid[96], grid[97], grid[113], grid[128], grid[129], grid[112]);
evolve8 e113 (grid_evolve[113], grid[96], grid[97], grid[98], grid[112], grid[114], grid[128], grid[129], grid[130], grid[113]);
evolve8 e114 (grid_evolve[114], grid[97], grid[98], grid[99], grid[113], grid[115], grid[129], grid[130], grid[131], grid[114]);
evolve8 e115 (grid_evolve[115], grid[98], grid[99], grid[100], grid[114], grid[116], grid[130], grid[131], grid[132], grid[115]);
evolve8 e116 (grid_evolve[116], grid[99], grid[100], grid[101], grid[115], grid[117], grid[131], grid[132], grid[133], grid[116]);
evolve8 e117 (grid_evolve[117], grid[100], grid[101], grid[102], grid[116], grid[118], grid[132], grid[133], grid[134], grid[117]);
evolve8 e118 (grid_evolve[118], grid[101], grid[102], grid[103], grid[117], grid[119], grid[133], grid[134], grid[135], grid[118]);
evolve8 e119 (grid_evolve[119], grid[102], grid[103], grid[104], grid[118], grid[120], grid[134], grid[135], grid[136], grid[119]);
evolve8 e120 (grid_evolve[120], grid[103], grid[104], grid[105], grid[119], grid[121], grid[135], grid[136], grid[137], grid[120]);
evolve8 e121 (grid_evolve[121], grid[104], grid[105], grid[106], grid[120], grid[122], grid[136], grid[137], grid[138], grid[121]);
evolve8 e122 (grid_evolve[122], grid[105], grid[106], grid[107], grid[121], grid[123], grid[137], grid[138], grid[139], grid[122]);
evolve8 e123 (grid_evolve[123], grid[106], grid[107], grid[108], grid[122], grid[124], grid[138], grid[139], grid[140], grid[123]);
evolve8 e124 (grid_evolve[124], grid[107], grid[108], grid[109], grid[123], grid[125], grid[139], grid[140], grid[141], grid[124]);
evolve8 e125 (grid_evolve[125], grid[108], grid[109], grid[110], grid[124], grid[126], grid[140], grid[141], grid[142], grid[125]);
evolve8 e126 (grid_evolve[126], grid[109], grid[110], grid[111], grid[125], grid[127], grid[141], grid[142], grid[143], grid[126]);
evolve5 e127 (grid_evolve[127], grid[110], grid[111], grid[126], grid[142], grid[143], grid[127]);

//row 9
evolve5 e128 (grid_evolve[128], grid[112], grid[113], grid[129], grid[144], grid[145], grid[128]);
evolve8 e129 (grid_evolve[129], grid[112], grid[113], grid[114], grid[128], grid[130], grid[144], grid[145], grid[146], grid[129]);
evolve8 e130 (grid_evolve[130], grid[113], grid[114], grid[115], grid[129], grid[131], grid[145], grid[146], grid[147], grid[130]);
evolve8 e131 (grid_evolve[131], grid[114], grid[115], grid[116], grid[130], grid[132], grid[146], grid[147], grid[148], grid[131]);
evolve8 e132 (grid_evolve[132], grid[115], grid[116], grid[117], grid[131], grid[133], grid[147], grid[148], grid[149], grid[132]);
evolve8 e133 (grid_evolve[133], grid[116], grid[117], grid[118], grid[132], grid[134], grid[148], grid[149], grid[150], grid[133]);
evolve8 e134 (grid_evolve[134], grid[117], grid[118], grid[119], grid[133], grid[135], grid[149], grid[150], grid[151], grid[134]);
evolve8 e135 (grid_evolve[135], grid[118], grid[119], grid[120], grid[134], grid[136], grid[150], grid[151], grid[152], grid[135]);
evolve8 e136 (grid_evolve[136], grid[119], grid[120], grid[121], grid[135], grid[137], grid[151], grid[152], grid[153], grid[136]);
evolve8 e137 (grid_evolve[137], grid[120], grid[121], grid[122], grid[136], grid[138], grid[152], grid[153], grid[154], grid[137]);
evolve8 e138 (grid_evolve[138], grid[121], grid[122], grid[123], grid[137], grid[139], grid[153], grid[154], grid[155], grid[138]);
evolve8 e139 (grid_evolve[139], grid[122], grid[123], grid[124], grid[138], grid[140], grid[154], grid[155], grid[156], grid[139]);
evolve8 e140 (grid_evolve[140], grid[123], grid[124], grid[125], grid[139], grid[141], grid[155], grid[156], grid[157], grid[140]);
evolve8 e141 (grid_evolve[141], grid[124], grid[125], grid[126], grid[140], grid[142], grid[156], grid[157], grid[158], grid[141]);
evolve8 e142 (grid_evolve[142], grid[125], grid[126], grid[127], grid[141], grid[143], grid[157], grid[158], grid[159], grid[142]);
evolve5 e143 (grid_evolve[143], grid[126], grid[127], grid[142], grid[158], grid[159], grid[143]);

//row 10
evolve5 e144 (grid_evolve[144], grid[128], grid[129], grid[145], grid[160], grid[161], grid[144]);
evolve8 e145 (grid_evolve[145], grid[128], grid[129], grid[130], grid[144], grid[146], grid[160], grid[161], grid[162], grid[145]);
evolve8 e146 (grid_evolve[146], grid[129], grid[130], grid[131], grid[145], grid[147], grid[161], grid[162], grid[163], grid[146]);
evolve8 e147 (grid_evolve[147], grid[130], grid[131], grid[132], grid[146], grid[148], grid[162], grid[163], grid[164], grid[147]);
evolve8 e148 (grid_evolve[148], grid[131], grid[132], grid[133], grid[147], grid[149], grid[163], grid[164], grid[165], grid[148]);
evolve8 e149 (grid_evolve[149], grid[132], grid[133], grid[134], grid[148], grid[150], grid[164], grid[165], grid[166], grid[149]);
evolve8 e150 (grid_evolve[150], grid[133], grid[134], grid[135], grid[149], grid[151], grid[165], grid[166], grid[167], grid[150]);
evolve8 e151 (grid_evolve[151], grid[134], grid[135], grid[136], grid[150], grid[152], grid[166], grid[167], grid[168], grid[151]);
evolve8 e152 (grid_evolve[152], grid[135], grid[136], grid[137], grid[151], grid[153], grid[167], grid[168], grid[169], grid[152]);
evolve8 e153 (grid_evolve[153], grid[136], grid[137], grid[138], grid[152], grid[154], grid[168], grid[169], grid[170], grid[153]);
evolve8 e154 (grid_evolve[154], grid[137], grid[138], grid[139], grid[153], grid[155], grid[169], grid[170], grid[171], grid[154]);
evolve8 e155 (grid_evolve[155], grid[138], grid[139], grid[140], grid[154], grid[156], grid[170], grid[171], grid[172], grid[155]);
evolve8 e156 (grid_evolve[156], grid[139], grid[140], grid[141], grid[155], grid[157], grid[171], grid[172], grid[173], grid[156]);
evolve8 e157 (grid_evolve[157], grid[140], grid[141], grid[142], grid[156], grid[158], grid[172], grid[173], grid[174], grid[157]);
evolve8 e158 (grid_evolve[158], grid[141], grid[142], grid[143], grid[157], grid[159], grid[173], grid[174], grid[175], grid[158]);
evolve5 e159 (grid_evolve[159], grid[142], grid[143], grid[158], grid[174], grid[175], grid[159]);

//row 11
evolve5 e160 (grid_evolve[160], grid[144], grid[145], grid[161], grid[176], grid[177], grid[160]);
evolve8 e161 (grid_evolve[161], grid[144], grid[145], grid[146], grid[160], grid[162], grid[176], grid[177], grid[178], grid[161]);
evolve8 e162 (grid_evolve[162], grid[145], grid[146], grid[147], grid[161], grid[163], grid[177], grid[178], grid[179], grid[162]);
evolve8 e163 (grid_evolve[163], grid[146], grid[147], grid[148], grid[162], grid[164], grid[178], grid[179], grid[180], grid[163]);
evolve8 e164 (grid_evolve[164], grid[147], grid[148], grid[149], grid[163], grid[165], grid[179], grid[180], grid[181], grid[164]);
evolve8 e165 (grid_evolve[165], grid[148], grid[149], grid[150], grid[164], grid[166], grid[180], grid[181], grid[182], grid[165]);
evolve8 e166 (grid_evolve[166], grid[149], grid[150], grid[151], grid[165], grid[167], grid[181], grid[182], grid[183], grid[166]);
evolve8 e167 (grid_evolve[167], grid[150], grid[151], grid[152], grid[166], grid[168], grid[182], grid[183], grid[184], grid[167]);
evolve8 e168 (grid_evolve[168], grid[151], grid[152], grid[153], grid[167], grid[169], grid[183], grid[184], grid[185], grid[168]);
evolve8 e169 (grid_evolve[169], grid[152], grid[153], grid[154], grid[168], grid[170], grid[184], grid[185], grid[186], grid[169]);
evolve8 e170 (grid_evolve[170], grid[153], grid[154], grid[155], grid[169], grid[171], grid[185], grid[186], grid[187], grid[170]);
evolve8 e171 (grid_evolve[171], grid[154], grid[155], grid[156], grid[170], grid[172], grid[186], grid[187], grid[188], grid[171]);
evolve8 e172 (grid_evolve[172], grid[155], grid[156], grid[157], grid[171], grid[173], grid[187], grid[188], grid[189], grid[172]);
evolve8 e173 (grid_evolve[173], grid[156], grid[157], grid[158], grid[172], grid[174], grid[188], grid[189], grid[190], grid[173]);
evolve8 e174 (grid_evolve[174], grid[157], grid[158], grid[159], grid[173], grid[175], grid[189], grid[190], grid[191], grid[174]);
evolve5 e175 (grid_evolve[175], grid[158], grid[159], grid[174], grid[190], grid[191], grid[175]);

//row 12
evolve5 e176 (grid_evolve[176], grid[160], grid[161], grid[177], grid[192], grid[193], grid[176]);
evolve8 e177 (grid_evolve[177], grid[160], grid[161], grid[162], grid[176], grid[178], grid[192], grid[193], grid[194], grid[177]);
evolve8 e178 (grid_evolve[178], grid[161], grid[162], grid[163], grid[177], grid[179], grid[193], grid[194], grid[195], grid[178]);
evolve8 e179 (grid_evolve[179], grid[162], grid[163], grid[164], grid[178], grid[180], grid[194], grid[195], grid[196], grid[179]);
evolve8 e180 (grid_evolve[180], grid[163], grid[164], grid[165], grid[179], grid[181], grid[195], grid[196], grid[197], grid[180]);
evolve8 e181 (grid_evolve[181], grid[164], grid[165], grid[166], grid[180], grid[182], grid[196], grid[197], grid[198], grid[181]);
evolve8 e182 (grid_evolve[182], grid[165], grid[166], grid[167], grid[181], grid[183], grid[197], grid[198], grid[199], grid[182]);
evolve8 e183 (grid_evolve[183], grid[166], grid[167], grid[168], grid[182], grid[184], grid[198], grid[199], grid[200], grid[183]);
evolve8 e184 (grid_evolve[184], grid[167], grid[168], grid[169], grid[183], grid[185], grid[199], grid[200], grid[201], grid[184]);
evolve8 e185 (grid_evolve[185], grid[168], grid[169], grid[170], grid[184], grid[186], grid[200], grid[201], grid[202], grid[185]);
evolve8 e186 (grid_evolve[186], grid[169], grid[170], grid[171], grid[185], grid[187], grid[201], grid[202], grid[203], grid[186]);
evolve8 e187 (grid_evolve[187], grid[170], grid[171], grid[172], grid[186], grid[188], grid[202], grid[203], grid[204], grid[187]);
evolve8 e188 (grid_evolve[188], grid[171], grid[172], grid[173], grid[187], grid[189], grid[203], grid[204], grid[205], grid[188]);
evolve8 e189 (grid_evolve[189], grid[172], grid[173], grid[174], grid[188], grid[190], grid[204], grid[205], grid[206], grid[189]);
evolve8 e190 (grid_evolve[190], grid[173], grid[174], grid[175], grid[189], grid[191], grid[205], grid[206], grid[207], grid[190]);
evolve5 e191 (grid_evolve[191], grid[174], grid[175], grid[190], grid[206], grid[207], grid[191]);

//row 13
evolve5 e192 (grid_evolve[192], grid[176], grid[177], grid[193], grid[208], grid[209], grid[192]);
evolve8 e193 (grid_evolve[193], grid[176], grid[177], grid[178], grid[192], grid[194], grid[208], grid[209], grid[210], grid[193]);
evolve8 e194 (grid_evolve[194], grid[177], grid[178], grid[179], grid[193], grid[195], grid[209], grid[210], grid[211], grid[194]);
evolve8 e195 (grid_evolve[195], grid[178], grid[179], grid[180], grid[194], grid[196], grid[210], grid[211], grid[212], grid[195]);
evolve8 e196 (grid_evolve[196], grid[179], grid[180], grid[181], grid[195], grid[197], grid[211], grid[212], grid[213], grid[196]);
evolve8 e197 (grid_evolve[197], grid[180], grid[181], grid[182], grid[196], grid[198], grid[212], grid[213], grid[214], grid[197]);
evolve8 e198 (grid_evolve[198], grid[181], grid[182], grid[183], grid[197], grid[199], grid[213], grid[214], grid[215], grid[198]);
evolve8 e199 (grid_evolve[199], grid[182], grid[183], grid[184], grid[198], grid[200], grid[214], grid[215], grid[216], grid[199]);
evolve8 e200 (grid_evolve[200], grid[183], grid[184], grid[185], grid[199], grid[201], grid[215], grid[216], grid[217], grid[200]);
evolve8 e201 (grid_evolve[201], grid[184], grid[185], grid[186], grid[200], grid[202], grid[216], grid[217], grid[218], grid[201]);
evolve8 e202 (grid_evolve[202], grid[185], grid[186], grid[187], grid[201], grid[203], grid[217], grid[218], grid[219], grid[202]);
evolve8 e203 (grid_evolve[203], grid[186], grid[187], grid[188], grid[202], grid[204], grid[218], grid[219], grid[220], grid[203]);
evolve8 e204 (grid_evolve[204], grid[187], grid[188], grid[189], grid[203], grid[205], grid[219], grid[220], grid[221], grid[204]);
evolve8 e205 (grid_evolve[205], grid[188], grid[189], grid[190], grid[204], grid[206], grid[220], grid[221], grid[222], grid[205]);
evolve8 e206 (grid_evolve[206], grid[189], grid[190], grid[191], grid[205], grid[207], grid[221], grid[222], grid[223], grid[206]);
evolve5 e207 (grid_evolve[207], grid[190], grid[191], grid[206], grid[222], grid[223], grid[207]);

//row 14
evolve5 e208 (grid_evolve[208], grid[192], grid[193], grid[209], grid[224], grid[225], grid[208]);
evolve8 e209 (grid_evolve[209], grid[192], grid[193], grid[194], grid[208], grid[210], grid[224], grid[225], grid[226], grid[209]);
evolve8 e210 (grid_evolve[210], grid[193], grid[194], grid[195], grid[209], grid[211], grid[225], grid[226], grid[227], grid[210]);
evolve8 e211 (grid_evolve[211], grid[194], grid[195], grid[196], grid[210], grid[212], grid[226], grid[227], grid[228], grid[211]);
evolve8 e212 (grid_evolve[212], grid[195], grid[196], grid[197], grid[211], grid[213], grid[227], grid[228], grid[229], grid[212]);
evolve8 e213 (grid_evolve[213], grid[196], grid[197], grid[198], grid[212], grid[214], grid[228], grid[229], grid[230], grid[213]);
evolve8 e214 (grid_evolve[214], grid[197], grid[198], grid[199], grid[213], grid[215], grid[229], grid[230], grid[231], grid[214]);
evolve8 e215 (grid_evolve[215], grid[198], grid[199], grid[200], grid[214], grid[216], grid[230], grid[231], grid[232], grid[215]);
evolve8 e216 (grid_evolve[216], grid[199], grid[200], grid[201], grid[215], grid[217], grid[231], grid[232], grid[233], grid[216]);
evolve8 e217 (grid_evolve[217], grid[200], grid[201], grid[202], grid[216], grid[218], grid[232], grid[233], grid[234], grid[217]);
evolve8 e218 (grid_evolve[218], grid[201], grid[202], grid[203], grid[217], grid[219], grid[233], grid[234], grid[235], grid[218]);
evolve8 e219 (grid_evolve[219], grid[202], grid[203], grid[204], grid[218], grid[220], grid[234], grid[235], grid[236], grid[219]);
evolve8 e220 (grid_evolve[220], grid[203], grid[204], grid[205], grid[219], grid[221], grid[235], grid[236], grid[237], grid[220]);
evolve8 e221 (grid_evolve[221], grid[204], grid[205], grid[206], grid[220], grid[222], grid[236], grid[237], grid[238], grid[221]);
evolve8 e222 (grid_evolve[222], grid[205], grid[206], grid[207], grid[221], grid[223], grid[237], grid[238], grid[239], grid[222]);
evolve5 e223 (grid_evolve[223], grid[206], grid[207], grid[222], grid[238], grid[239], grid[223]);

//row 15
evolve5 e224 (grid_evolve[224], grid[208], grid[209], grid[225], grid[240], grid[241], grid[224]);
evolve8 e225 (grid_evolve[225], grid[208], grid[209], grid[210], grid[224], grid[226], grid[240], grid[241], grid[242], grid[225]);
evolve8 e226 (grid_evolve[226], grid[209], grid[210], grid[211], grid[225], grid[227], grid[241], grid[242], grid[243], grid[226]);
evolve8 e227 (grid_evolve[227], grid[210], grid[211], grid[212], grid[226], grid[228], grid[242], grid[243], grid[244], grid[227]);
evolve8 e228 (grid_evolve[228], grid[211], grid[212], grid[213], grid[227], grid[229], grid[243], grid[244], grid[245], grid[228]);
evolve8 e229 (grid_evolve[229], grid[212], grid[213], grid[214], grid[228], grid[230], grid[244], grid[245], grid[246], grid[229]);
evolve8 e230 (grid_evolve[230], grid[213], grid[214], grid[215], grid[229], grid[231], grid[245], grid[246], grid[247], grid[230]);
evolve8 e231 (grid_evolve[231], grid[214], grid[215], grid[216], grid[230], grid[232], grid[246], grid[247], grid[248], grid[231]);
evolve8 e232 (grid_evolve[232], grid[215], grid[216], grid[217], grid[231], grid[233], grid[247], grid[248], grid[249], grid[232]);
evolve8 e233 (grid_evolve[233], grid[216], grid[217], grid[218], grid[232], grid[234], grid[248], grid[249], grid[250], grid[233]);
evolve8 e234 (grid_evolve[234], grid[217], grid[218], grid[219], grid[233], grid[235], grid[249], grid[250], grid[251], grid[234]);
evolve8 e235 (grid_evolve[235], grid[218], grid[219], grid[220], grid[234], grid[236], grid[250], grid[251], grid[252], grid[235]);
evolve8 e236 (grid_evolve[236], grid[219], grid[220], grid[221], grid[235], grid[237], grid[251], grid[252], grid[253], grid[236]);
evolve8 e237 (grid_evolve[237], grid[220], grid[221], grid[222], grid[236], grid[238], grid[252], grid[253], grid[254], grid[237]);
evolve8 e238 (grid_evolve[238], grid[221], grid[222], grid[223], grid[237], grid[239], grid[253], grid[254], grid[255], grid[238]);
evolve5 e239 (grid_evolve[239], grid[222], grid[223], grid[238], grid[254], grid[255], grid[239]);

//row 16
evolve3 e240 (grid_evolve[240], grid[224], grid[225], grid[241], grid[240]);
evolve5 e241 (grid_evolve[241], grid[224], grid[225], grid[226], grid[240], grid[242], grid[241]);
evolve5 e242 (grid_evolve[242], grid[225], grid[226], grid[227], grid[241], grid[243], grid[242]);
evolve5 e243 (grid_evolve[243], grid[226], grid[227], grid[228], grid[242], grid[244], grid[243]);
evolve5 e244 (grid_evolve[244], grid[227], grid[228], grid[229], grid[243], grid[245], grid[244]);
evolve5 e245 (grid_evolve[245], grid[228], grid[229], grid[230], grid[244], grid[246], grid[245]);
evolve5 e246 (grid_evolve[246], grid[229], grid[230], grid[231], grid[245], grid[247], grid[246]);
evolve5 e247 (grid_evolve[247], grid[230], grid[231], grid[232], grid[246], grid[248], grid[247]);
evolve5 e248 (grid_evolve[248], grid[231], grid[232], grid[233], grid[247], grid[249], grid[248]);
evolve5 e249 (grid_evolve[249], grid[232], grid[233], grid[234], grid[248], grid[250], grid[249]);
evolve5 e250 (grid_evolve[250], grid[233], grid[234], grid[235], grid[249], grid[251], grid[250]);
evolve5 e251 (grid_evolve[251], grid[234], grid[235], grid[236], grid[250], grid[252], grid[251]);
evolve5 e252 (grid_evolve[252], grid[235], grid[236], grid[237], grid[251], grid[253], grid[252]);
evolve5 e253 (grid_evolve[253], grid[236], grid[237], grid[238], grid[252], grid[254], grid[253]);
evolve5 e254 (grid_evolve[254], grid[237], grid[238], grid[239], grid[253], grid[255], grid[254]);
evolve3 e255 (grid_evolve[255], grid[238], grid[239], grid[254], grid[255]);
 
endmodule // top


module evolve3 (next_state, vector1, vector2, vector3, current_state);
	
   input logic  vector1;
   input logic  vector2;
   input logic  vector3;
   input logic  current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve3

module evolve5 (next_state, vector1, vector2, vector3, 
		vector4, vector5, current_state);
   
   input logic     vector1;
   input logic 	 vector2;
   input logic 	 vector3;
   input logic 	 vector4;
   input logic 	 vector5;
   input logic 	 current_state;
   output logic    next_state;
   
   logic [3:0] 	 sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + vector5;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve5


module evolve8 (next_state, vector1, vector2, vector3, 
		vector4, vector5, vector6, 
		vector7, vector8, current_state);
   
   input logic 	vector1;
   input logic 	vector2;
   input logic 	vector3;
   input logic 	vector4;
   input logic 	vector5;
	
   input logic 	vector6;
   input logic 	vector7;
   input logic 	vector8;
   input logic 	current_state;
   output logic   next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + 
		vector5 + vector6 + vector7 + vector8;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve8


module rules (pop_count, current_state, next_state);
   
   input logic [3:0] pop_count;
   input logic 	     current_state;
   output logic      next_state;
   
   assign next_state = (pop_count == 2 & current_state) | pop_count == 3;
   
endmodule // rules