/*
 
 Conway's Game of Life modeled in SVerilog
 
 */
module datapath (clk, mux2out, initial_seed, run, reset);
input logic clk;
input logic [575:0]  initial_seed;
input logic          reset;
input logic          run;
output logic [575:0] mux2out;

logic [575:0] 	grid;
logic [575:0]   grid_evolve, ffout;
logic start_or_cont;
logic en;

   evolve efga (grid, grid_evolve);
   fsm f1 (clk, run, reset, start_or_cont, en);
   mux2 #(576)m1 (ffout, initial_seed, start_or_cont, grid);
   mux2 #(576)m2 (ffout, initial_seed, reset, mux2out);
   flopen #(576)flop1 (clk, en, grid_evolve, ffout);

endmodule

module fsm (clk, run, reset, start_or_cont, en);

input logic clk;
input logic          reset;
input logic          run;
output logic         start_or_cont;
output logic         en; 

typedef enum 	logic [1:0] {S0, S1, S2, S3} statetype;
   statetype state, nextstate;
   
   // state register
   always_ff @(posedge clk, posedge reset)
     if (reset) state <= S0;
     else state <= nextstate;
   
   // next state logic
   always_comb
     case (state)
       S0: begin 
         if(run) begin
          nextstate <= S1;
          start_or_cont = 1'b1;
          en = 1'b1;
         end
         else begin 
          nextstate <= S0;
          start_or_cont = 1'b1;
          en = 1'b1;
         end
       end

       S1: begin
         if(run) begin 
          nextstate <= S1;
          start_or_cont = 1'b0;
          en = 1'b1;
         end
         else if(run == 0) begin 
          nextstate <= S2;
          start_or_cont = 1'b0;
          en = 1'b1;
         end
         else begin 
          nextstate <= S0;
          start_or_cont = 1'b1;
          en = 1'b1;
         end
       end

       S2: begin
         if(run) begin 
          nextstate <= S1;
         end
         else if(run == 0) begin 
          nextstate <= S2;
          start_or_cont = 1'b0;
          en = 1'b0;
         end
         else begin
          nextstate <= S0;
         end
       end

       S3: begin
         nextstate <= S0;
       end
     endcase

endmodule

module mux2 #(parameter WIDTH = 8) (
  input  logic [WIDTH-1:0] d0, d1, 
  input  logic             s, 
  output logic [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule

`timescale 1ns / 1ps
module flopen #(parameter WIDTH = 8) (
  input  logic             clk, en,
  input  logic [WIDTH-1:0] d, 
  output logic [WIDTH-1:0] q);

  always_ff @(posedge clk)
    if (en) q <= #1 d;
    else q <= q;
endmodule

module evolve (grid, grid_evolve);
input logic [575:0] 	grid;
output logic [575:0] 	grid_evolve;
//row 1  
evolve3 e0 (grid_evolve[0], grid[1], grid[24], grid[25], grid[0]);
evolve5 e1 (grid_evolve[1], grid[0], grid[2], grid[24], grid[25], grid[26], grid[1]);
evolve5 e2 (grid_evolve[2], grid[1], grid[3], grid[25], grid[26], grid[27], grid[2]);
evolve5 e3 (grid_evolve[3], grid[2], grid[4], grid[26], grid[27], grid[28], grid[3]);
evolve5 e4 (grid_evolve[4], grid[3], grid[5], grid[27], grid[28], grid[29], grid[4]);
evolve5 e5 (grid_evolve[5], grid[4], grid[6], grid[28], grid[29], grid[30], grid[5]);
evolve5 e6 (grid_evolve[6], grid[5], grid[7], grid[29], grid[30], grid[31], grid[6]);
evolve5 e7 (grid_evolve[7], grid[6], grid[8], grid[30], grid[31], grid[32], grid[7]);
evolve5 e8 (grid_evolve[8], grid[7], grid[9], grid[31], grid[32], grid[33], grid[8]);
evolve5 e9 (grid_evolve[9], grid[8], grid[10], grid[32], grid[33], grid[34], grid[9]);
evolve5 e10 (grid_evolve[10], grid[9], grid[11], grid[33], grid[34], grid[35], grid[10]);
evolve5 e11 (grid_evolve[11], grid[10], grid[12], grid[34], grid[35], grid[36], grid[11]);
evolve5 e12 (grid_evolve[12], grid[11], grid[13], grid[35], grid[36], grid[37], grid[12]);
evolve5 e13 (grid_evolve[13], grid[12], grid[14], grid[36], grid[37], grid[38], grid[13]);
evolve5 e14 (grid_evolve[14], grid[13], grid[15], grid[37], grid[38], grid[39], grid[14]);
evolve5 e15 (grid_evolve[15], grid[14], grid[16], grid[38], grid[39], grid[40], grid[15]);
evolve5 e16 (grid_evolve[16], grid[15], grid[17], grid[39], grid[40], grid[41], grid[16]);
evolve5 e17 (grid_evolve[17], grid[16], grid[18], grid[40], grid[41], grid[42], grid[17]);
evolve5 e18 (grid_evolve[18], grid[17], grid[19], grid[41], grid[42], grid[43], grid[18]);
evolve5 e19 (grid_evolve[19], grid[18], grid[20], grid[42], grid[43], grid[44], grid[19]);
evolve5 e20 (grid_evolve[20], grid[19], grid[21], grid[43], grid[44], grid[45], grid[20]);
evolve5 e21 (grid_evolve[21], grid[20], grid[22], grid[44], grid[45], grid[46], grid[21]);
evolve5 e22 (grid_evolve[22], grid[21], grid[23], grid[45], grid[46], grid[47], grid[22]);
evolve3 e23 (grid_evolve[23], grid[22], grid[46], grid[47], grid[23]);

evolve5 e24 (grid_evolve[24], grid[0], grid[1], grid[25], grid[48], grid[49], grid[24]);
evolve8 e25 (grid_evolve[25], grid[0], grid[1], grid[2], grid[24], grid[26], grid[48], grid[49], grid[50], grid[25]);
evolve8 e26 (grid_evolve[26], grid[1], grid[2], grid[3], grid[25], grid[27], grid[49], grid[50], grid[51], grid[26]);
evolve8 e27 (grid_evolve[27], grid[2], grid[3], grid[4], grid[26], grid[28], grid[50], grid[51], grid[52], grid[27]);
evolve8 e28 (grid_evolve[28], grid[3], grid[4], grid[5], grid[27], grid[29], grid[51], grid[52], grid[53], grid[28]);
evolve8 e29 (grid_evolve[29], grid[4], grid[5], grid[6], grid[28], grid[30], grid[52], grid[53], grid[54], grid[29]);
evolve8 e30 (grid_evolve[30], grid[5], grid[6], grid[7], grid[29], grid[31], grid[53], grid[54], grid[55], grid[30]);
evolve8 e31 (grid_evolve[31], grid[6], grid[7], grid[8], grid[30], grid[32], grid[54], grid[55], grid[56], grid[31]);
evolve8 e32 (grid_evolve[32], grid[7], grid[8], grid[9], grid[31], grid[33], grid[55], grid[56], grid[57], grid[32]);
evolve8 e33 (grid_evolve[33], grid[8], grid[9], grid[10], grid[32], grid[34], grid[56], grid[57], grid[58], grid[33]);
evolve8 e34 (grid_evolve[34], grid[9], grid[10], grid[11], grid[33], grid[35], grid[57], grid[58], grid[59], grid[34]);
evolve8 e35 (grid_evolve[35], grid[10], grid[11], grid[12], grid[34], grid[36], grid[58], grid[59], grid[60], grid[35]);
evolve8 e36 (grid_evolve[36], grid[11], grid[12], grid[13], grid[35], grid[37], grid[59], grid[60], grid[61], grid[36]);
evolve8 e37 (grid_evolve[37], grid[12], grid[13], grid[14], grid[36], grid[38], grid[60], grid[61], grid[62], grid[37]);
evolve8 e38 (grid_evolve[38], grid[13], grid[14], grid[15], grid[37], grid[39], grid[61], grid[62], grid[63], grid[38]);
evolve8 e39 (grid_evolve[39], grid[14], grid[15], grid[16], grid[38], grid[40], grid[62], grid[63], grid[64], grid[39]);
evolve8 e40 (grid_evolve[40], grid[15], grid[16], grid[17], grid[39], grid[41], grid[63], grid[64], grid[65], grid[40]);
evolve8 e41 (grid_evolve[41], grid[16], grid[17], grid[18], grid[40], grid[42], grid[64], grid[65], grid[66], grid[41]);
evolve8 e42 (grid_evolve[42], grid[17], grid[18], grid[19], grid[41], grid[43], grid[65], grid[66], grid[67], grid[42]);
evolve8 e43 (grid_evolve[43], grid[18], grid[19], grid[20], grid[42], grid[44], grid[66], grid[67], grid[68], grid[43]);
evolve8 e44 (grid_evolve[44], grid[19], grid[20], grid[21], grid[43], grid[45], grid[67], grid[68], grid[69], grid[44]);
evolve8 e45 (grid_evolve[45], grid[20], grid[21], grid[22], grid[44], grid[46], grid[68], grid[69], grid[70], grid[45]);
evolve8 e46 (grid_evolve[46], grid[21], grid[22], grid[23], grid[45], grid[47], grid[69], grid[70], grid[71], grid[46]);
evolve5 e47 (grid_evolve[47], grid[22], grid[23], grid[46], grid[70], grid[71], grid[47]);
evolve5 e48 (grid_evolve[48], grid[24], grid[25], grid[49], grid[72], grid[73], grid[48]);
evolve8 e49 (grid_evolve[49], grid[24], grid[25], grid[26], grid[48], grid[50], grid[72], grid[73], grid[74], grid[49]);
evolve8 e50 (grid_evolve[50], grid[25], grid[26], grid[27], grid[49], grid[51], grid[73], grid[74], grid[75], grid[50]);
evolve8 e51 (grid_evolve[51], grid[26], grid[27], grid[28], grid[50], grid[52], grid[74], grid[75], grid[76], grid[51]);
evolve8 e52 (grid_evolve[52], grid[27], grid[28], grid[29], grid[51], grid[53], grid[75], grid[76], grid[77], grid[52]);
evolve8 e53 (grid_evolve[53], grid[28], grid[29], grid[30], grid[52], grid[54], grid[76], grid[77], grid[78], grid[53]);
evolve8 e54 (grid_evolve[54], grid[29], grid[30], grid[31], grid[53], grid[55], grid[77], grid[78], grid[79], grid[54]);
evolve8 e55 (grid_evolve[55], grid[30], grid[31], grid[32], grid[54], grid[56], grid[78], grid[79], grid[80], grid[55]);
evolve8 e56 (grid_evolve[56], grid[31], grid[32], grid[33], grid[55], grid[57], grid[79], grid[80], grid[81], grid[56]);
evolve8 e57 (grid_evolve[57], grid[32], grid[33], grid[34], grid[56], grid[58], grid[80], grid[81], grid[82], grid[57]);
evolve8 e58 (grid_evolve[58], grid[33], grid[34], grid[35], grid[57], grid[59], grid[81], grid[82], grid[83], grid[58]);
evolve8 e59 (grid_evolve[59], grid[34], grid[35], grid[36], grid[58], grid[60], grid[82], grid[83], grid[84], grid[59]);
evolve8 e60 (grid_evolve[60], grid[35], grid[36], grid[37], grid[59], grid[61], grid[83], grid[84], grid[85], grid[60]);
evolve8 e61 (grid_evolve[61], grid[36], grid[37], grid[38], grid[60], grid[62], grid[84], grid[85], grid[86], grid[61]);
evolve8 e62 (grid_evolve[62], grid[37], grid[38], grid[39], grid[61], grid[63], grid[85], grid[86], grid[87], grid[62]);
evolve8 e63 (grid_evolve[63], grid[38], grid[39], grid[40], grid[62], grid[64], grid[86], grid[87], grid[88], grid[63]);
evolve8 e64 (grid_evolve[64], grid[39], grid[40], grid[41], grid[63], grid[65], grid[87], grid[88], grid[89], grid[64]);
evolve8 e65 (grid_evolve[65], grid[40], grid[41], grid[42], grid[64], grid[66], grid[88], grid[89], grid[90], grid[65]);
evolve8 e66 (grid_evolve[66], grid[41], grid[42], grid[43], grid[65], grid[67], grid[89], grid[90], grid[91], grid[66]);
evolve8 e67 (grid_evolve[67], grid[42], grid[43], grid[44], grid[66], grid[68], grid[90], grid[91], grid[92], grid[67]);
evolve8 e68 (grid_evolve[68], grid[43], grid[44], grid[45], grid[67], grid[69], grid[91], grid[92], grid[93], grid[68]);
evolve8 e69 (grid_evolve[69], grid[44], grid[45], grid[46], grid[68], grid[70], grid[92], grid[93], grid[94], grid[69]);
evolve8 e70 (grid_evolve[70], grid[45], grid[46], grid[47], grid[69], grid[71], grid[93], grid[94], grid[95], grid[70]);
evolve5 e71 (grid_evolve[71], grid[46], grid[47], grid[70], grid[94], grid[95], grid[71]);

evolve5 e72 (grid_evolve[72], grid[48], grid[49], grid[73], grid[96], grid[97], grid[72]);
evolve8 e73 (grid_evolve[73], grid[48], grid[49], grid[50], grid[72], grid[74], grid[96], grid[97], grid[98], grid[73]);
evolve8 e74 (grid_evolve[74], grid[49], grid[50], grid[51], grid[73], grid[75], grid[97], grid[98], grid[99], grid[74]);
evolve8 e75 (grid_evolve[75], grid[50], grid[51], grid[52], grid[74], grid[76], grid[98], grid[99], grid[100], grid[75]);
evolve8 e76 (grid_evolve[76], grid[51], grid[52], grid[53], grid[75], grid[77], grid[99], grid[100], grid[101], grid[76]);
evolve8 e77 (grid_evolve[77], grid[52], grid[53], grid[54], grid[76], grid[78], grid[100], grid[101], grid[102], grid[77]);
evolve8 e78 (grid_evolve[78], grid[53], grid[54], grid[55], grid[77], grid[79], grid[101], grid[102], grid[103], grid[78]);
evolve8 e79 (grid_evolve[79], grid[54], grid[55], grid[56], grid[78], grid[80], grid[102], grid[103], grid[104], grid[79]);
evolve8 e80 (grid_evolve[80], grid[55], grid[56], grid[57], grid[79], grid[81], grid[103], grid[104], grid[105], grid[80]);
evolve8 e81 (grid_evolve[81], grid[56], grid[57], grid[58], grid[80], grid[82], grid[104], grid[105], grid[106], grid[81]);
evolve8 e82 (grid_evolve[82], grid[57], grid[58], grid[59], grid[81], grid[83], grid[105], grid[106], grid[107], grid[82]);
evolve8 e83 (grid_evolve[83], grid[58], grid[59], grid[60], grid[82], grid[84], grid[106], grid[107], grid[108], grid[83]);
evolve8 e84 (grid_evolve[84], grid[59], grid[60], grid[61], grid[83], grid[85], grid[107], grid[108], grid[109], grid[84]);
evolve8 e85 (grid_evolve[85], grid[60], grid[61], grid[62], grid[84], grid[86], grid[108], grid[109], grid[110], grid[85]);
evolve8 e86 (grid_evolve[86], grid[61], grid[62], grid[63], grid[85], grid[87], grid[109], grid[110], grid[111], grid[86]);
evolve8 e87 (grid_evolve[87], grid[62], grid[63], grid[64], grid[86], grid[88], grid[110], grid[111], grid[112], grid[87]);
evolve8 e88 (grid_evolve[88], grid[63], grid[64], grid[65], grid[87], grid[89], grid[111], grid[112], grid[113], grid[88]);
evolve8 e89 (grid_evolve[89], grid[64], grid[65], grid[66], grid[88], grid[90], grid[112], grid[113], grid[114], grid[89]);
evolve8 e90 (grid_evolve[90], grid[65], grid[66], grid[67], grid[89], grid[91], grid[113], grid[114], grid[115], grid[90]);
evolve8 e91 (grid_evolve[91], grid[66], grid[67], grid[68], grid[90], grid[92], grid[114], grid[115], grid[116], grid[91]);
evolve8 e92 (grid_evolve[92], grid[67], grid[68], grid[69], grid[91], grid[93], grid[115], grid[116], grid[117], grid[92]);
evolve8 e93 (grid_evolve[93], grid[68], grid[69], grid[70], grid[92], grid[94], grid[116], grid[117], grid[118], grid[93]);
evolve8 e94 (grid_evolve[94], grid[69], grid[70], grid[71], grid[93], grid[95], grid[117], grid[118], grid[119], grid[94]);
evolve5 e95 (grid_evolve[95], grid[70], grid[71], grid[94], grid[118], grid[119], grid[95]);

evolve5 e96 (grid_evolve[96], grid[72], grid[73], grid[97], grid[120], grid[121], grid[96]);
evolve8 e97 (grid_evolve[97], grid[72], grid[73], grid[74], grid[96], grid[98], grid[120], grid[121], grid[122], grid[97]);
evolve8 e98 (grid_evolve[98], grid[73], grid[74], grid[75], grid[97], grid[99], grid[121], grid[122], grid[123], grid[98]);
evolve8 e99 (grid_evolve[99], grid[74], grid[75], grid[76], grid[98], grid[100], grid[122], grid[123], grid[124], grid[99]);
evolve8 e100 (grid_evolve[100], grid[75], grid[76], grid[77], grid[99], grid[101], grid[123], grid[124], grid[125], grid[100]);
evolve8 e101 (grid_evolve[101], grid[76], grid[77], grid[78], grid[100], grid[102], grid[124], grid[125], grid[126], grid[101]);
evolve8 e102 (grid_evolve[102], grid[77], grid[78], grid[79], grid[101], grid[103], grid[125], grid[126], grid[127], grid[102]);
evolve8 e103 (grid_evolve[103], grid[78], grid[79], grid[80], grid[102], grid[104], grid[126], grid[127], grid[128], grid[103]);
evolve8 e104 (grid_evolve[104], grid[79], grid[80], grid[81], grid[103], grid[105], grid[127], grid[128], grid[129], grid[104]);
evolve8 e105 (grid_evolve[105], grid[80], grid[81], grid[82], grid[104], grid[106], grid[128], grid[129], grid[130], grid[105]);
evolve8 e106 (grid_evolve[106], grid[81], grid[82], grid[83], grid[105], grid[107], grid[129], grid[130], grid[131], grid[106]);
evolve8 e107 (grid_evolve[107], grid[82], grid[83], grid[84], grid[106], grid[108], grid[130], grid[131], grid[132], grid[107]);
evolve8 e108 (grid_evolve[108], grid[83], grid[84], grid[85], grid[107], grid[109], grid[131], grid[132], grid[133], grid[108]);
evolve8 e109 (grid_evolve[109], grid[84], grid[85], grid[86], grid[108], grid[110], grid[132], grid[133], grid[134], grid[109]);
evolve8 e110 (grid_evolve[110], grid[85], grid[86], grid[87], grid[109], grid[111], grid[133], grid[134], grid[135], grid[110]);
evolve8 e111 (grid_evolve[111], grid[86], grid[87], grid[88], grid[110], grid[112], grid[134], grid[135], grid[136], grid[111]);
evolve8 e112 (grid_evolve[112], grid[87], grid[88], grid[89], grid[111], grid[113], grid[135], grid[136], grid[137], grid[112]);
evolve8 e113 (grid_evolve[113], grid[88], grid[89], grid[90], grid[112], grid[114], grid[136], grid[137], grid[138], grid[113]);
evolve8 e114 (grid_evolve[114], grid[89], grid[90], grid[91], grid[113], grid[115], grid[137], grid[138], grid[139], grid[114]);
evolve8 e115 (grid_evolve[115], grid[90], grid[91], grid[92], grid[114], grid[116], grid[138], grid[139], grid[140], grid[115]);
evolve8 e116 (grid_evolve[116], grid[91], grid[92], grid[93], grid[115], grid[117], grid[139], grid[140], grid[141], grid[116]);
evolve8 e117 (grid_evolve[117], grid[92], grid[93], grid[94], grid[116], grid[118], grid[140], grid[141], grid[142], grid[117]);
evolve8 e118 (grid_evolve[118], grid[93], grid[94], grid[95], grid[117], grid[119], grid[141], grid[142], grid[143], grid[118]);
evolve5 e119 (grid_evolve[119], grid[94], grid[95], grid[118], grid[142], grid[143], grid[119]);

evolve5 e120 (grid_evolve[120], grid[96], grid[97], grid[121], grid[144], grid[145], grid[120]);
evolve8 e121 (grid_evolve[121], grid[96], grid[97], grid[98], grid[120], grid[122], grid[144], grid[145], grid[146], grid[121]);
evolve8 e122 (grid_evolve[122], grid[97], grid[98], grid[99], grid[121], grid[123], grid[145], grid[146], grid[147], grid[122]);
evolve8 e123 (grid_evolve[123], grid[98], grid[99], grid[100], grid[122], grid[124], grid[146], grid[147], grid[148], grid[123]);
evolve8 e124 (grid_evolve[124], grid[99], grid[100], grid[101], grid[123], grid[125], grid[147], grid[148], grid[149], grid[124]);
evolve8 e125 (grid_evolve[125], grid[100], grid[101], grid[102], grid[124], grid[126], grid[148], grid[149], grid[150], grid[125]);
evolve8 e126 (grid_evolve[126], grid[101], grid[102], grid[103], grid[125], grid[127], grid[149], grid[150], grid[151], grid[126]);
evolve8 e127 (grid_evolve[127], grid[102], grid[103], grid[104], grid[126], grid[128], grid[150], grid[151], grid[152], grid[127]);
evolve8 e128 (grid_evolve[128], grid[103], grid[104], grid[105], grid[127], grid[129], grid[151], grid[152], grid[153], grid[128]);
evolve8 e129 (grid_evolve[129], grid[104], grid[105], grid[106], grid[128], grid[130], grid[152], grid[153], grid[154], grid[129]);
evolve8 e130 (grid_evolve[130], grid[105], grid[106], grid[107], grid[129], grid[131], grid[153], grid[154], grid[155], grid[130]);
evolve8 e131 (grid_evolve[131], grid[106], grid[107], grid[108], grid[130], grid[132], grid[154], grid[155], grid[156], grid[131]);
evolve8 e132 (grid_evolve[132], grid[107], grid[108], grid[109], grid[131], grid[133], grid[155], grid[156], grid[157], grid[132]);
evolve8 e133 (grid_evolve[133], grid[108], grid[109], grid[110], grid[132], grid[134], grid[156], grid[157], grid[158], grid[133]);
evolve8 e134 (grid_evolve[134], grid[109], grid[110], grid[111], grid[133], grid[135], grid[157], grid[158], grid[159], grid[134]);
evolve8 e135 (grid_evolve[135], grid[110], grid[111], grid[112], grid[134], grid[136], grid[158], grid[159], grid[160], grid[135]);
evolve8 e136 (grid_evolve[136], grid[111], grid[112], grid[113], grid[135], grid[137], grid[159], grid[160], grid[161], grid[136]);
evolve8 e137 (grid_evolve[137], grid[112], grid[113], grid[114], grid[136], grid[138], grid[160], grid[161], grid[162], grid[137]);
evolve8 e138 (grid_evolve[138], grid[113], grid[114], grid[115], grid[137], grid[139], grid[161], grid[162], grid[163], grid[138]);
evolve8 e139 (grid_evolve[139], grid[114], grid[115], grid[116], grid[138], grid[140], grid[162], grid[163], grid[164], grid[139]);
evolve8 e140 (grid_evolve[140], grid[115], grid[116], grid[117], grid[139], grid[141], grid[163], grid[164], grid[165], grid[140]);
evolve8 e141 (grid_evolve[141], grid[116], grid[117], grid[118], grid[140], grid[142], grid[164], grid[165], grid[166], grid[141]);
evolve8 e142 (grid_evolve[142], grid[117], grid[118], grid[119], grid[141], grid[143], grid[165], grid[166], grid[167], grid[142]);
evolve5 e143 (grid_evolve[143], grid[118], grid[119], grid[142], grid[166], grid[167], grid[143]);

evolve5 e144 (grid_evolve[144], grid[120], grid[121], grid[145], grid[168], grid[169], grid[144]);
evolve8 e145 (grid_evolve[145], grid[120], grid[121], grid[122], grid[144], grid[146], grid[168], grid[169], grid[170], grid[145]);
evolve8 e146 (grid_evolve[146], grid[121], grid[122], grid[123], grid[145], grid[147], grid[169], grid[170], grid[171], grid[146]);
evolve8 e147 (grid_evolve[147], grid[122], grid[123], grid[124], grid[146], grid[148], grid[170], grid[171], grid[172], grid[147]);
evolve8 e148 (grid_evolve[148], grid[123], grid[124], grid[125], grid[147], grid[149], grid[171], grid[172], grid[173], grid[148]);
evolve8 e149 (grid_evolve[149], grid[124], grid[125], grid[126], grid[148], grid[150], grid[172], grid[173], grid[174], grid[149]);
evolve8 e150 (grid_evolve[150], grid[125], grid[126], grid[127], grid[149], grid[151], grid[173], grid[174], grid[175], grid[150]);
evolve8 e151 (grid_evolve[151], grid[126], grid[127], grid[128], grid[150], grid[152], grid[174], grid[175], grid[176], grid[151]);
evolve8 e152 (grid_evolve[152], grid[127], grid[128], grid[129], grid[151], grid[153], grid[175], grid[176], grid[177], grid[152]);
evolve8 e153 (grid_evolve[153], grid[128], grid[129], grid[130], grid[152], grid[154], grid[176], grid[177], grid[178], grid[153]);
evolve8 e154 (grid_evolve[154], grid[129], grid[130], grid[131], grid[153], grid[155], grid[177], grid[178], grid[179], grid[154]);
evolve8 e155 (grid_evolve[155], grid[130], grid[131], grid[132], grid[154], grid[156], grid[178], grid[179], grid[180], grid[155]);
evolve8 e156 (grid_evolve[156], grid[131], grid[132], grid[133], grid[155], grid[157], grid[179], grid[180], grid[181], grid[156]);
evolve8 e157 (grid_evolve[157], grid[132], grid[133], grid[134], grid[156], grid[158], grid[180], grid[181], grid[182], grid[157]);
evolve8 e158 (grid_evolve[158], grid[133], grid[134], grid[135], grid[157], grid[159], grid[181], grid[182], grid[183], grid[158]);
evolve8 e159 (grid_evolve[159], grid[134], grid[135], grid[136], grid[158], grid[160], grid[182], grid[183], grid[184], grid[159]);
evolve8 e160 (grid_evolve[160], grid[135], grid[136], grid[137], grid[159], grid[161], grid[183], grid[184], grid[185], grid[160]);
evolve8 e161 (grid_evolve[161], grid[136], grid[137], grid[138], grid[160], grid[162], grid[184], grid[185], grid[186], grid[161]);
evolve8 e162 (grid_evolve[162], grid[137], grid[138], grid[139], grid[161], grid[163], grid[185], grid[186], grid[187], grid[162]);
evolve8 e163 (grid_evolve[163], grid[138], grid[139], grid[140], grid[162], grid[164], grid[186], grid[187], grid[188], grid[163]);
evolve8 e164 (grid_evolve[164], grid[139], grid[140], grid[141], grid[163], grid[165], grid[187], grid[188], grid[189], grid[164]);
evolve8 e165 (grid_evolve[165], grid[140], grid[141], grid[142], grid[164], grid[166], grid[188], grid[189], grid[190], grid[165]);
evolve8 e166 (grid_evolve[166], grid[141], grid[142], grid[143], grid[165], grid[167], grid[189], grid[190], grid[191], grid[166]);
evolve5 e167 (grid_evolve[167], grid[142], grid[143], grid[166], grid[190], grid[191], grid[167]);

evolve5 e168 (grid_evolve[168], grid[144], grid[145], grid[169], grid[192], grid[193], grid[168]);
evolve8 e169 (grid_evolve[169], grid[144], grid[145], grid[146], grid[168], grid[170], grid[192], grid[193], grid[194], grid[169]);
evolve8 e170 (grid_evolve[170], grid[145], grid[146], grid[147], grid[169], grid[171], grid[193], grid[194], grid[195], grid[170]);
evolve8 e171 (grid_evolve[171], grid[146], grid[147], grid[148], grid[170], grid[172], grid[194], grid[195], grid[196], grid[171]);
evolve8 e172 (grid_evolve[172], grid[147], grid[148], grid[149], grid[171], grid[173], grid[195], grid[196], grid[197], grid[172]);
evolve8 e173 (grid_evolve[173], grid[148], grid[149], grid[150], grid[172], grid[174], grid[196], grid[197], grid[198], grid[173]);
evolve8 e174 (grid_evolve[174], grid[149], grid[150], grid[151], grid[173], grid[175], grid[197], grid[198], grid[199], grid[174]);
evolve8 e175 (grid_evolve[175], grid[150], grid[151], grid[152], grid[174], grid[176], grid[198], grid[199], grid[200], grid[175]);
evolve8 e176 (grid_evolve[176], grid[151], grid[152], grid[153], grid[175], grid[177], grid[199], grid[200], grid[201], grid[176]);
evolve8 e177 (grid_evolve[177], grid[152], grid[153], grid[154], grid[176], grid[178], grid[200], grid[201], grid[202], grid[177]);
evolve8 e178 (grid_evolve[178], grid[153], grid[154], grid[155], grid[177], grid[179], grid[201], grid[202], grid[203], grid[178]);
evolve8 e179 (grid_evolve[179], grid[154], grid[155], grid[156], grid[178], grid[180], grid[202], grid[203], grid[204], grid[179]);
evolve8 e180 (grid_evolve[180], grid[155], grid[156], grid[157], grid[179], grid[181], grid[203], grid[204], grid[205], grid[180]);
evolve8 e181 (grid_evolve[181], grid[156], grid[157], grid[158], grid[180], grid[182], grid[204], grid[205], grid[206], grid[181]);
evolve8 e182 (grid_evolve[182], grid[157], grid[158], grid[159], grid[181], grid[183], grid[205], grid[206], grid[207], grid[182]);
evolve8 e183 (grid_evolve[183], grid[158], grid[159], grid[160], grid[182], grid[184], grid[206], grid[207], grid[208], grid[183]);
evolve8 e184 (grid_evolve[184], grid[159], grid[160], grid[161], grid[183], grid[185], grid[207], grid[208], grid[209], grid[184]);
evolve8 e185 (grid_evolve[185], grid[160], grid[161], grid[162], grid[184], grid[186], grid[208], grid[209], grid[210], grid[185]);
evolve8 e186 (grid_evolve[186], grid[161], grid[162], grid[163], grid[185], grid[187], grid[209], grid[210], grid[211], grid[186]);
evolve8 e187 (grid_evolve[187], grid[162], grid[163], grid[164], grid[186], grid[188], grid[210], grid[211], grid[212], grid[187]);
evolve8 e188 (grid_evolve[188], grid[163], grid[164], grid[165], grid[187], grid[189], grid[211], grid[212], grid[213], grid[188]);
evolve8 e189 (grid_evolve[189], grid[164], grid[165], grid[166], grid[188], grid[190], grid[212], grid[213], grid[214], grid[189]);
evolve8 e190 (grid_evolve[190], grid[165], grid[166], grid[167], grid[189], grid[191], grid[213], grid[214], grid[215], grid[190]);
evolve5 e191 (grid_evolve[191], grid[166], grid[167], grid[190], grid[214], grid[215], grid[191]);

evolve5 e192 (grid_evolve[192], grid[168], grid[169], grid[193], grid[216], grid[217], grid[192]);
evolve8 e193 (grid_evolve[193], grid[168], grid[169], grid[170], grid[192], grid[194], grid[216], grid[217], grid[218], grid[193]);
evolve8 e194 (grid_evolve[194], grid[169], grid[170], grid[171], grid[193], grid[195], grid[217], grid[218], grid[219], grid[194]);
evolve8 e195 (grid_evolve[195], grid[170], grid[171], grid[172], grid[194], grid[196], grid[218], grid[219], grid[220], grid[195]);
evolve8 e196 (grid_evolve[196], grid[171], grid[172], grid[173], grid[195], grid[197], grid[219], grid[220], grid[221], grid[196]);
evolve8 e197 (grid_evolve[197], grid[172], grid[173], grid[174], grid[196], grid[198], grid[220], grid[221], grid[222], grid[197]);
evolve8 e198 (grid_evolve[198], grid[173], grid[174], grid[175], grid[197], grid[199], grid[221], grid[222], grid[223], grid[198]);
evolve8 e199 (grid_evolve[199], grid[174], grid[175], grid[176], grid[198], grid[200], grid[222], grid[223], grid[224], grid[199]);
evolve8 e200 (grid_evolve[200], grid[175], grid[176], grid[177], grid[199], grid[201], grid[223], grid[224], grid[225], grid[200]);
evolve8 e201 (grid_evolve[201], grid[176], grid[177], grid[178], grid[200], grid[202], grid[224], grid[225], grid[226], grid[201]);
evolve8 e202 (grid_evolve[202], grid[177], grid[178], grid[179], grid[201], grid[203], grid[225], grid[226], grid[227], grid[202]);
evolve8 e203 (grid_evolve[203], grid[178], grid[179], grid[180], grid[202], grid[204], grid[226], grid[227], grid[228], grid[203]);
evolve8 e204 (grid_evolve[204], grid[179], grid[180], grid[181], grid[203], grid[205], grid[227], grid[228], grid[229], grid[204]);
evolve8 e205 (grid_evolve[205], grid[180], grid[181], grid[182], grid[204], grid[206], grid[228], grid[229], grid[230], grid[205]);
evolve8 e206 (grid_evolve[206], grid[181], grid[182], grid[183], grid[205], grid[207], grid[229], grid[230], grid[231], grid[206]);
evolve8 e207 (grid_evolve[207], grid[182], grid[183], grid[184], grid[206], grid[208], grid[230], grid[231], grid[232], grid[207]);
evolve8 e208 (grid_evolve[208], grid[183], grid[184], grid[185], grid[207], grid[209], grid[231], grid[232], grid[233], grid[208]);
evolve8 e209 (grid_evolve[209], grid[184], grid[185], grid[186], grid[208], grid[210], grid[232], grid[233], grid[234], grid[209]);
evolve8 e210 (grid_evolve[210], grid[185], grid[186], grid[187], grid[209], grid[211], grid[233], grid[234], grid[235], grid[210]);
evolve8 e211 (grid_evolve[211], grid[186], grid[187], grid[188], grid[210], grid[212], grid[234], grid[235], grid[236], grid[211]);
evolve8 e212 (grid_evolve[212], grid[187], grid[188], grid[189], grid[211], grid[213], grid[235], grid[236], grid[237], grid[212]);
evolve8 e213 (grid_evolve[213], grid[188], grid[189], grid[190], grid[212], grid[214], grid[236], grid[237], grid[238], grid[213]);
evolve8 e214 (grid_evolve[214], grid[189], grid[190], grid[191], grid[213], grid[215], grid[237], grid[238], grid[239], grid[214]);
evolve5 e215 (grid_evolve[215], grid[190], grid[191], grid[214], grid[238], grid[239], grid[215]);

evolve5 e216 (grid_evolve[216], grid[192], grid[193], grid[217], grid[240], grid[241], grid[216]);
evolve8 e217 (grid_evolve[217], grid[192], grid[193], grid[194], grid[216], grid[218], grid[240], grid[241], grid[242], grid[217]);
evolve8 e218 (grid_evolve[218], grid[193], grid[194], grid[195], grid[217], grid[219], grid[241], grid[242], grid[243], grid[218]);
evolve8 e219 (grid_evolve[219], grid[194], grid[195], grid[196], grid[218], grid[220], grid[242], grid[243], grid[244], grid[219]);
evolve8 e220 (grid_evolve[220], grid[195], grid[196], grid[197], grid[219], grid[221], grid[243], grid[244], grid[245], grid[220]);
evolve8 e221 (grid_evolve[221], grid[196], grid[197], grid[198], grid[220], grid[222], grid[244], grid[245], grid[246], grid[221]);
evolve8 e222 (grid_evolve[222], grid[197], grid[198], grid[199], grid[221], grid[223], grid[245], grid[246], grid[247], grid[222]);
evolve8 e223 (grid_evolve[223], grid[198], grid[199], grid[200], grid[222], grid[224], grid[246], grid[247], grid[248], grid[223]);
evolve8 e224 (grid_evolve[224], grid[199], grid[200], grid[201], grid[223], grid[225], grid[247], grid[248], grid[249], grid[224]);
evolve8 e225 (grid_evolve[225], grid[200], grid[201], grid[202], grid[224], grid[226], grid[248], grid[249], grid[250], grid[225]);
evolve8 e226 (grid_evolve[226], grid[201], grid[202], grid[203], grid[225], grid[227], grid[249], grid[250], grid[251], grid[226]);
evolve8 e227 (grid_evolve[227], grid[202], grid[203], grid[204], grid[226], grid[228], grid[250], grid[251], grid[252], grid[227]);
evolve8 e228 (grid_evolve[228], grid[203], grid[204], grid[205], grid[227], grid[229], grid[251], grid[252], grid[253], grid[228]);
evolve8 e229 (grid_evolve[229], grid[204], grid[205], grid[206], grid[228], grid[230], grid[252], grid[253], grid[254], grid[229]);
evolve8 e230 (grid_evolve[230], grid[205], grid[206], grid[207], grid[229], grid[231], grid[253], grid[254], grid[255], grid[230]);
evolve8 e231 (grid_evolve[231], grid[206], grid[207], grid[208], grid[230], grid[232], grid[254], grid[255], grid[256], grid[231]);
evolve8 e232 (grid_evolve[232], grid[207], grid[208], grid[209], grid[231], grid[233], grid[255], grid[256], grid[257], grid[232]);
evolve8 e233 (grid_evolve[233], grid[208], grid[209], grid[210], grid[232], grid[234], grid[256], grid[257], grid[258], grid[233]);
evolve8 e234 (grid_evolve[234], grid[209], grid[210], grid[211], grid[233], grid[235], grid[257], grid[258], grid[259], grid[234]);
evolve8 e235 (grid_evolve[235], grid[210], grid[211], grid[212], grid[234], grid[236], grid[258], grid[259], grid[260], grid[235]);
evolve8 e236 (grid_evolve[236], grid[211], grid[212], grid[213], grid[235], grid[237], grid[259], grid[260], grid[261], grid[236]);
evolve8 e237 (grid_evolve[237], grid[212], grid[213], grid[214], grid[236], grid[238], grid[260], grid[261], grid[262], grid[237]);
evolve8 e238 (grid_evolve[238], grid[213], grid[214], grid[215], grid[237], grid[239], grid[261], grid[262], grid[263], grid[238]);
evolve5 e239 (grid_evolve[239], grid[214], grid[215], grid[238], grid[262], grid[263], grid[239]);

evolve5 e240 (grid_evolve[240], grid[216], grid[217], grid[241], grid[264], grid[265], grid[240]);
evolve8 e241 (grid_evolve[241], grid[216], grid[217], grid[218], grid[240], grid[242], grid[264], grid[265], grid[266], grid[241]);
evolve8 e242 (grid_evolve[242], grid[217], grid[218], grid[219], grid[241], grid[243], grid[265], grid[266], grid[267], grid[242]);
evolve8 e243 (grid_evolve[243], grid[218], grid[219], grid[220], grid[242], grid[244], grid[266], grid[267], grid[268], grid[243]);
evolve8 e244 (grid_evolve[244], grid[219], grid[220], grid[221], grid[243], grid[245], grid[267], grid[268], grid[269], grid[244]);
evolve8 e245 (grid_evolve[245], grid[220], grid[221], grid[222], grid[244], grid[246], grid[268], grid[269], grid[270], grid[245]);
evolve8 e246 (grid_evolve[246], grid[221], grid[222], grid[223], grid[245], grid[247], grid[269], grid[270], grid[271], grid[246]);
evolve8 e247 (grid_evolve[247], grid[222], grid[223], grid[224], grid[246], grid[248], grid[270], grid[271], grid[272], grid[247]);
evolve8 e248 (grid_evolve[248], grid[223], grid[224], grid[225], grid[247], grid[249], grid[271], grid[272], grid[273], grid[248]);
evolve8 e249 (grid_evolve[249], grid[224], grid[225], grid[226], grid[248], grid[250], grid[272], grid[273], grid[274], grid[249]);
evolve8 e250 (grid_evolve[250], grid[225], grid[226], grid[227], grid[249], grid[251], grid[273], grid[274], grid[275], grid[250]);
evolve8 e251 (grid_evolve[251], grid[226], grid[227], grid[228], grid[250], grid[252], grid[274], grid[275], grid[276], grid[251]);
evolve8 e252 (grid_evolve[252], grid[227], grid[228], grid[229], grid[251], grid[253], grid[275], grid[276], grid[277], grid[252]);
evolve8 e253 (grid_evolve[253], grid[228], grid[229], grid[230], grid[252], grid[254], grid[276], grid[277], grid[278], grid[253]);
evolve8 e254 (grid_evolve[254], grid[229], grid[230], grid[231], grid[253], grid[255], grid[277], grid[278], grid[279], grid[254]);
evolve8 e255 (grid_evolve[255], grid[230], grid[231], grid[232], grid[254], grid[256], grid[278], grid[279], grid[280], grid[255]);
evolve8 e256 (grid_evolve[256], grid[231], grid[232], grid[233], grid[255], grid[257], grid[279], grid[280], grid[281], grid[256]);
evolve8 e257 (grid_evolve[257], grid[232], grid[233], grid[234], grid[256], grid[258], grid[280], grid[281], grid[282], grid[257]);
evolve8 e258 (grid_evolve[258], grid[233], grid[234], grid[235], grid[257], grid[259], grid[281], grid[282], grid[283], grid[258]);
evolve8 e259 (grid_evolve[259], grid[234], grid[235], grid[236], grid[258], grid[260], grid[282], grid[283], grid[284], grid[259]);
evolve8 e260 (grid_evolve[260], grid[235], grid[236], grid[237], grid[259], grid[261], grid[283], grid[284], grid[285], grid[260]);
evolve8 e261 (grid_evolve[261], grid[236], grid[237], grid[238], grid[260], grid[262], grid[284], grid[285], grid[286], grid[261]);
evolve8 e262 (grid_evolve[262], grid[237], grid[238], grid[239], grid[261], grid[263], grid[285], grid[286], grid[287], grid[262]);
evolve5 e263 (grid_evolve[263], grid[238], grid[239], grid[262], grid[286], grid[287], grid[263]);

evolve5 e264 (grid_evolve[264], grid[240], grid[241], grid[265], grid[288], grid[289], grid[264]);
evolve8 e265 (grid_evolve[265], grid[240], grid[241], grid[242], grid[264], grid[266], grid[288], grid[289], grid[290], grid[265]);
evolve8 e266 (grid_evolve[266], grid[241], grid[242], grid[243], grid[265], grid[267], grid[289], grid[290], grid[291], grid[266]);
evolve8 e267 (grid_evolve[267], grid[242], grid[243], grid[244], grid[266], grid[268], grid[290], grid[291], grid[292], grid[267]);
evolve8 e268 (grid_evolve[268], grid[243], grid[244], grid[245], grid[267], grid[269], grid[291], grid[292], grid[293], grid[268]);
evolve8 e269 (grid_evolve[269], grid[244], grid[245], grid[246], grid[268], grid[270], grid[292], grid[293], grid[294], grid[269]);
evolve8 e270 (grid_evolve[270], grid[245], grid[246], grid[247], grid[269], grid[271], grid[293], grid[294], grid[295], grid[270]);
evolve8 e271 (grid_evolve[271], grid[246], grid[247], grid[248], grid[270], grid[272], grid[294], grid[295], grid[296], grid[271]);
evolve8 e272 (grid_evolve[272], grid[247], grid[248], grid[249], grid[271], grid[273], grid[295], grid[296], grid[297], grid[272]);
evolve8 e273 (grid_evolve[273], grid[248], grid[249], grid[250], grid[272], grid[274], grid[296], grid[297], grid[298], grid[273]);
evolve8 e274 (grid_evolve[274], grid[249], grid[250], grid[251], grid[273], grid[275], grid[297], grid[298], grid[299], grid[274]);
evolve8 e275 (grid_evolve[275], grid[250], grid[251], grid[252], grid[274], grid[276], grid[298], grid[299], grid[300], grid[275]);
evolve8 e276 (grid_evolve[276], grid[251], grid[252], grid[253], grid[275], grid[277], grid[299], grid[300], grid[301], grid[276]);
evolve8 e277 (grid_evolve[277], grid[252], grid[253], grid[254], grid[276], grid[278], grid[300], grid[301], grid[302], grid[277]);
evolve8 e278 (grid_evolve[278], grid[253], grid[254], grid[255], grid[277], grid[279], grid[301], grid[302], grid[303], grid[278]);
evolve8 e279 (grid_evolve[279], grid[254], grid[255], grid[256], grid[278], grid[280], grid[302], grid[303], grid[304], grid[279]);
evolve8 e280 (grid_evolve[280], grid[255], grid[256], grid[257], grid[279], grid[281], grid[303], grid[304], grid[305], grid[280]);
evolve8 e281 (grid_evolve[281], grid[256], grid[257], grid[258], grid[280], grid[282], grid[304], grid[305], grid[306], grid[281]);
evolve8 e282 (grid_evolve[282], grid[257], grid[258], grid[259], grid[281], grid[283], grid[305], grid[306], grid[307], grid[282]);
evolve8 e283 (grid_evolve[283], grid[258], grid[259], grid[260], grid[282], grid[284], grid[306], grid[307], grid[308], grid[283]);
evolve8 e284 (grid_evolve[284], grid[259], grid[260], grid[261], grid[283], grid[285], grid[307], grid[308], grid[309], grid[284]);
evolve8 e285 (grid_evolve[285], grid[260], grid[261], grid[262], grid[284], grid[286], grid[308], grid[309], grid[310], grid[285]);
evolve8 e286 (grid_evolve[286], grid[261], grid[262], grid[263], grid[285], grid[287], grid[309], grid[310], grid[311], grid[286]);
evolve5 e287 (grid_evolve[287], grid[262], grid[263], grid[286], grid[310], grid[311], grid[287]);

evolve5 e288 (grid_evolve[288], grid[264], grid[265], grid[289], grid[312], grid[313], grid[288]);
evolve8 e289 (grid_evolve[289], grid[264], grid[265], grid[266], grid[288], grid[290], grid[312], grid[313], grid[314], grid[289]);
evolve8 e290 (grid_evolve[290], grid[265], grid[266], grid[267], grid[289], grid[291], grid[313], grid[314], grid[315], grid[290]);
evolve8 e291 (grid_evolve[291], grid[266], grid[267], grid[268], grid[290], grid[292], grid[314], grid[315], grid[316], grid[291]);
evolve8 e292 (grid_evolve[292], grid[267], grid[268], grid[269], grid[291], grid[293], grid[315], grid[316], grid[317], grid[292]);
evolve8 e293 (grid_evolve[293], grid[268], grid[269], grid[270], grid[292], grid[294], grid[316], grid[317], grid[318], grid[293]);
evolve8 e294 (grid_evolve[294], grid[269], grid[270], grid[271], grid[293], grid[295], grid[317], grid[318], grid[319], grid[294]);
evolve8 e295 (grid_evolve[295], grid[270], grid[271], grid[272], grid[294], grid[296], grid[318], grid[319], grid[320], grid[295]);
evolve8 e296 (grid_evolve[296], grid[271], grid[272], grid[273], grid[295], grid[297], grid[319], grid[320], grid[321], grid[296]);
evolve8 e297 (grid_evolve[297], grid[272], grid[273], grid[274], grid[296], grid[298], grid[320], grid[321], grid[322], grid[297]);
evolve8 e298 (grid_evolve[298], grid[273], grid[274], grid[275], grid[297], grid[299], grid[321], grid[322], grid[323], grid[298]);
evolve8 e299 (grid_evolve[299], grid[274], grid[275], grid[276], grid[298], grid[300], grid[322], grid[323], grid[324], grid[299]);
evolve8 e300 (grid_evolve[300], grid[275], grid[276], grid[277], grid[299], grid[301], grid[323], grid[324], grid[325], grid[300]);
evolve8 e301 (grid_evolve[301], grid[276], grid[277], grid[278], grid[300], grid[302], grid[324], grid[325], grid[326], grid[301]);
evolve8 e302 (grid_evolve[302], grid[277], grid[278], grid[279], grid[301], grid[303], grid[325], grid[326], grid[327], grid[302]);
evolve8 e303 (grid_evolve[303], grid[278], grid[279], grid[280], grid[302], grid[304], grid[326], grid[327], grid[328], grid[303]);
evolve8 e304 (grid_evolve[304], grid[279], grid[280], grid[281], grid[303], grid[305], grid[327], grid[328], grid[329], grid[304]);
evolve8 e305 (grid_evolve[305], grid[280], grid[281], grid[282], grid[304], grid[306], grid[328], grid[329], grid[330], grid[305]);
evolve8 e306 (grid_evolve[306], grid[281], grid[282], grid[283], grid[305], grid[307], grid[329], grid[330], grid[331], grid[306]);
evolve8 e307 (grid_evolve[307], grid[282], grid[283], grid[284], grid[306], grid[308], grid[330], grid[331], grid[332], grid[307]);
evolve8 e308 (grid_evolve[308], grid[283], grid[284], grid[285], grid[307], grid[309], grid[331], grid[332], grid[333], grid[308]);
evolve8 e309 (grid_evolve[309], grid[284], grid[285], grid[286], grid[308], grid[310], grid[332], grid[333], grid[334], grid[309]);
evolve8 e310 (grid_evolve[310], grid[285], grid[286], grid[287], grid[309], grid[311], grid[333], grid[334], grid[335], grid[310]);
evolve5 e311 (grid_evolve[311], grid[286], grid[287], grid[310], grid[334], grid[335], grid[311]);

evolve5 e312 (grid_evolve[312], grid[288], grid[289], grid[313], grid[336], grid[337], grid[312]);
evolve8 e313 (grid_evolve[313], grid[288], grid[289], grid[290], grid[312], grid[314], grid[336], grid[337], grid[338], grid[313]);
evolve8 e314 (grid_evolve[314], grid[289], grid[290], grid[291], grid[313], grid[315], grid[337], grid[338], grid[339], grid[314]);
evolve8 e315 (grid_evolve[315], grid[290], grid[291], grid[292], grid[314], grid[316], grid[338], grid[339], grid[340], grid[315]);
evolve8 e316 (grid_evolve[316], grid[291], grid[292], grid[293], grid[315], grid[317], grid[339], grid[340], grid[341], grid[316]);
evolve8 e317 (grid_evolve[317], grid[292], grid[293], grid[294], grid[316], grid[318], grid[340], grid[341], grid[342], grid[317]);
evolve8 e318 (grid_evolve[318], grid[293], grid[294], grid[295], grid[317], grid[319], grid[341], grid[342], grid[343], grid[318]);
evolve8 e319 (grid_evolve[319], grid[294], grid[295], grid[296], grid[318], grid[320], grid[342], grid[343], grid[344], grid[319]);
evolve8 e320 (grid_evolve[320], grid[295], grid[296], grid[297], grid[319], grid[321], grid[343], grid[344], grid[345], grid[320]);
evolve8 e321 (grid_evolve[321], grid[296], grid[297], grid[298], grid[320], grid[322], grid[344], grid[345], grid[346], grid[321]);
evolve8 e322 (grid_evolve[322], grid[297], grid[298], grid[299], grid[321], grid[323], grid[345], grid[346], grid[347], grid[322]);
evolve8 e323 (grid_evolve[323], grid[298], grid[299], grid[300], grid[322], grid[324], grid[346], grid[347], grid[348], grid[323]);
evolve8 e324 (grid_evolve[324], grid[299], grid[300], grid[301], grid[323], grid[325], grid[347], grid[348], grid[349], grid[324]);
evolve8 e325 (grid_evolve[325], grid[300], grid[301], grid[302], grid[324], grid[326], grid[348], grid[349], grid[350], grid[325]);
evolve8 e326 (grid_evolve[326], grid[301], grid[302], grid[303], grid[325], grid[327], grid[349], grid[350], grid[351], grid[326]);
evolve8 e327 (grid_evolve[327], grid[302], grid[303], grid[304], grid[326], grid[328], grid[350], grid[351], grid[352], grid[327]);
evolve8 e328 (grid_evolve[328], grid[303], grid[304], grid[305], grid[327], grid[329], grid[351], grid[352], grid[353], grid[328]);
evolve8 e329 (grid_evolve[329], grid[304], grid[305], grid[306], grid[328], grid[330], grid[352], grid[353], grid[354], grid[329]);
evolve8 e330 (grid_evolve[330], grid[305], grid[306], grid[307], grid[329], grid[331], grid[353], grid[354], grid[355], grid[330]);
evolve8 e331 (grid_evolve[331], grid[306], grid[307], grid[308], grid[330], grid[332], grid[354], grid[355], grid[356], grid[331]);
evolve8 e332 (grid_evolve[332], grid[307], grid[308], grid[309], grid[331], grid[333], grid[355], grid[356], grid[357], grid[332]);
evolve8 e333 (grid_evolve[333], grid[308], grid[309], grid[310], grid[332], grid[334], grid[356], grid[357], grid[358], grid[333]);
evolve8 e334 (grid_evolve[334], grid[309], grid[310], grid[311], grid[333], grid[335], grid[357], grid[358], grid[359], grid[334]);
evolve5 e335 (grid_evolve[335], grid[310], grid[311], grid[334], grid[358], grid[359], grid[335]);

evolve5 e336 (grid_evolve[336], grid[312], grid[313], grid[337], grid[360], grid[361], grid[336]);
evolve8 e337 (grid_evolve[337], grid[312], grid[313], grid[314], grid[336], grid[338], grid[360], grid[361], grid[362], grid[337]);
evolve8 e338 (grid_evolve[338], grid[313], grid[314], grid[315], grid[337], grid[339], grid[361], grid[362], grid[363], grid[338]);
evolve8 e339 (grid_evolve[339], grid[314], grid[315], grid[316], grid[338], grid[340], grid[362], grid[363], grid[364], grid[339]);
evolve8 e340 (grid_evolve[340], grid[315], grid[316], grid[317], grid[339], grid[341], grid[363], grid[364], grid[365], grid[340]);
evolve8 e341 (grid_evolve[341], grid[316], grid[317], grid[318], grid[340], grid[342], grid[364], grid[365], grid[366], grid[341]);
evolve8 e342 (grid_evolve[342], grid[317], grid[318], grid[319], grid[341], grid[343], grid[365], grid[366], grid[367], grid[342]);
evolve8 e343 (grid_evolve[343], grid[318], grid[319], grid[320], grid[342], grid[344], grid[366], grid[367], grid[368], grid[343]);
evolve8 e344 (grid_evolve[344], grid[319], grid[320], grid[321], grid[343], grid[345], grid[367], grid[368], grid[369], grid[344]);
evolve8 e345 (grid_evolve[345], grid[320], grid[321], grid[322], grid[344], grid[346], grid[368], grid[369], grid[370], grid[345]);
evolve8 e346 (grid_evolve[346], grid[321], grid[322], grid[323], grid[345], grid[347], grid[369], grid[370], grid[371], grid[346]);
evolve8 e347 (grid_evolve[347], grid[322], grid[323], grid[324], grid[346], grid[348], grid[370], grid[371], grid[372], grid[347]);
evolve8 e348 (grid_evolve[348], grid[323], grid[324], grid[325], grid[347], grid[349], grid[371], grid[372], grid[373], grid[348]);
evolve8 e349 (grid_evolve[349], grid[324], grid[325], grid[326], grid[348], grid[350], grid[372], grid[373], grid[374], grid[349]);
evolve8 e350 (grid_evolve[350], grid[325], grid[326], grid[327], grid[349], grid[351], grid[373], grid[374], grid[375], grid[350]);
evolve8 e351 (grid_evolve[351], grid[326], grid[327], grid[328], grid[350], grid[352], grid[374], grid[375], grid[376], grid[351]);
evolve8 e352 (grid_evolve[352], grid[327], grid[328], grid[329], grid[351], grid[353], grid[375], grid[376], grid[377], grid[352]);
evolve8 e353 (grid_evolve[353], grid[328], grid[329], grid[330], grid[352], grid[354], grid[376], grid[377], grid[378], grid[353]);
evolve8 e354 (grid_evolve[354], grid[329], grid[330], grid[331], grid[353], grid[355], grid[377], grid[378], grid[379], grid[354]);
evolve8 e355 (grid_evolve[355], grid[330], grid[331], grid[332], grid[354], grid[356], grid[378], grid[379], grid[380], grid[355]);
evolve8 e356 (grid_evolve[356], grid[331], grid[332], grid[333], grid[355], grid[357], grid[379], grid[380], grid[381], grid[356]);
evolve8 e357 (grid_evolve[357], grid[332], grid[333], grid[334], grid[356], grid[358], grid[380], grid[381], grid[382], grid[357]);
evolve8 e358 (grid_evolve[358], grid[333], grid[334], grid[335], grid[357], grid[359], grid[381], grid[382], grid[383], grid[358]);
evolve5 e359 (grid_evolve[359], grid[334], grid[335], grid[358], grid[382], grid[383], grid[359]);

evolve5 e360 (grid_evolve[360], grid[336], grid[337], grid[361], grid[384], grid[385], grid[360]);
evolve8 e361 (grid_evolve[361], grid[336], grid[337], grid[338], grid[360], grid[362], grid[384], grid[385], grid[386], grid[361]);
evolve8 e362 (grid_evolve[362], grid[337], grid[338], grid[339], grid[361], grid[363], grid[385], grid[386], grid[387], grid[362]);
evolve8 e363 (grid_evolve[363], grid[338], grid[339], grid[340], grid[362], grid[364], grid[386], grid[387], grid[388], grid[363]);
evolve8 e364 (grid_evolve[364], grid[339], grid[340], grid[341], grid[363], grid[365], grid[387], grid[388], grid[389], grid[364]);
evolve8 e365 (grid_evolve[365], grid[340], grid[341], grid[342], grid[364], grid[366], grid[388], grid[389], grid[390], grid[365]);
evolve8 e366 (grid_evolve[366], grid[341], grid[342], grid[343], grid[365], grid[367], grid[389], grid[390], grid[391], grid[366]);
evolve8 e367 (grid_evolve[367], grid[342], grid[343], grid[344], grid[366], grid[368], grid[390], grid[391], grid[392], grid[367]);
evolve8 e368 (grid_evolve[368], grid[343], grid[344], grid[345], grid[367], grid[369], grid[391], grid[392], grid[393], grid[368]);
evolve8 e369 (grid_evolve[369], grid[344], grid[345], grid[346], grid[368], grid[370], grid[392], grid[393], grid[394], grid[369]);
evolve8 e370 (grid_evolve[370], grid[345], grid[346], grid[347], grid[369], grid[371], grid[393], grid[394], grid[395], grid[370]);
evolve8 e371 (grid_evolve[371], grid[346], grid[347], grid[348], grid[370], grid[372], grid[394], grid[395], grid[396], grid[371]);
evolve8 e372 (grid_evolve[372], grid[347], grid[348], grid[349], grid[371], grid[373], grid[395], grid[396], grid[397], grid[372]);
evolve8 e373 (grid_evolve[373], grid[348], grid[349], grid[350], grid[372], grid[374], grid[396], grid[397], grid[398], grid[373]);
evolve8 e374 (grid_evolve[374], grid[349], grid[350], grid[351], grid[373], grid[375], grid[397], grid[398], grid[399], grid[374]);
evolve8 e375 (grid_evolve[375], grid[350], grid[351], grid[352], grid[374], grid[376], grid[398], grid[399], grid[400], grid[375]);
evolve8 e376 (grid_evolve[376], grid[351], grid[352], grid[353], grid[375], grid[377], grid[399], grid[400], grid[401], grid[376]);
evolve8 e377 (grid_evolve[377], grid[352], grid[353], grid[354], grid[376], grid[378], grid[400], grid[401], grid[402], grid[377]);
evolve8 e378 (grid_evolve[378], grid[353], grid[354], grid[355], grid[377], grid[379], grid[401], grid[402], grid[403], grid[378]);
evolve8 e379 (grid_evolve[379], grid[354], grid[355], grid[356], grid[378], grid[380], grid[402], grid[403], grid[404], grid[379]);
evolve8 e380 (grid_evolve[380], grid[355], grid[356], grid[357], grid[379], grid[381], grid[403], grid[404], grid[405], grid[380]);
evolve8 e381 (grid_evolve[381], grid[356], grid[357], grid[358], grid[380], grid[382], grid[404], grid[405], grid[406], grid[381]);
evolve8 e382 (grid_evolve[382], grid[357], grid[358], grid[359], grid[381], grid[383], grid[405], grid[406], grid[407], grid[382]);
evolve5 e383 (grid_evolve[383], grid[358], grid[359], grid[382], grid[406], grid[407], grid[383]);

evolve5 e384 (grid_evolve[384], grid[360], grid[361], grid[385], grid[408], grid[409], grid[384]);
evolve8 e385 (grid_evolve[385], grid[360], grid[361], grid[362], grid[384], grid[386], grid[408], grid[409], grid[410], grid[385]);
evolve8 e386 (grid_evolve[386], grid[361], grid[362], grid[363], grid[385], grid[387], grid[409], grid[410], grid[411], grid[386]);
evolve8 e387 (grid_evolve[387], grid[362], grid[363], grid[364], grid[386], grid[388], grid[410], grid[411], grid[412], grid[387]);
evolve8 e388 (grid_evolve[388], grid[363], grid[364], grid[365], grid[387], grid[389], grid[411], grid[412], grid[413], grid[388]);
evolve8 e389 (grid_evolve[389], grid[364], grid[365], grid[366], grid[388], grid[390], grid[412], grid[413], grid[414], grid[389]);
evolve8 e390 (grid_evolve[390], grid[365], grid[366], grid[367], grid[389], grid[391], grid[413], grid[414], grid[415], grid[390]);
evolve8 e391 (grid_evolve[391], grid[366], grid[367], grid[368], grid[390], grid[392], grid[414], grid[415], grid[416], grid[391]);
evolve8 e392 (grid_evolve[392], grid[367], grid[368], grid[369], grid[391], grid[393], grid[415], grid[416], grid[417], grid[392]);
evolve8 e393 (grid_evolve[393], grid[368], grid[369], grid[370], grid[392], grid[394], grid[416], grid[417], grid[418], grid[393]);
evolve8 e394 (grid_evolve[394], grid[369], grid[370], grid[371], grid[393], grid[395], grid[417], grid[418], grid[419], grid[394]);
evolve8 e395 (grid_evolve[395], grid[370], grid[371], grid[372], grid[394], grid[396], grid[418], grid[419], grid[420], grid[395]);
evolve8 e396 (grid_evolve[396], grid[371], grid[372], grid[373], grid[395], grid[397], grid[419], grid[420], grid[421], grid[396]);
evolve8 e397 (grid_evolve[397], grid[372], grid[373], grid[374], grid[396], grid[398], grid[420], grid[421], grid[422], grid[397]);
evolve8 e398 (grid_evolve[398], grid[373], grid[374], grid[375], grid[397], grid[399], grid[421], grid[422], grid[423], grid[398]);
evolve8 e399 (grid_evolve[399], grid[374], grid[375], grid[376], grid[398], grid[400], grid[422], grid[423], grid[424], grid[399]);
evolve8 e400 (grid_evolve[400], grid[375], grid[376], grid[377], grid[399], grid[401], grid[423], grid[424], grid[425], grid[400]);
evolve8 e401 (grid_evolve[401], grid[376], grid[377], grid[378], grid[400], grid[402], grid[424], grid[425], grid[426], grid[401]);
evolve8 e402 (grid_evolve[402], grid[377], grid[378], grid[379], grid[401], grid[403], grid[425], grid[426], grid[427], grid[402]);
evolve8 e403 (grid_evolve[403], grid[378], grid[379], grid[380], grid[402], grid[404], grid[426], grid[427], grid[428], grid[403]);
evolve8 e404 (grid_evolve[404], grid[379], grid[380], grid[381], grid[403], grid[405], grid[427], grid[428], grid[429], grid[404]);
evolve8 e405 (grid_evolve[405], grid[380], grid[381], grid[382], grid[404], grid[406], grid[428], grid[429], grid[430], grid[405]);
evolve8 e406 (grid_evolve[406], grid[381], grid[382], grid[383], grid[405], grid[407], grid[429], grid[430], grid[431], grid[406]);
evolve5 e407 (grid_evolve[407], grid[382], grid[383], grid[406], grid[430], grid[431], grid[407]);

evolve5 e408 (grid_evolve[408], grid[384], grid[385], grid[409], grid[432], grid[433], grid[408]);
evolve8 e409 (grid_evolve[409], grid[384], grid[385], grid[386], grid[408], grid[410], grid[432], grid[433], grid[434], grid[409]);
evolve8 e410 (grid_evolve[410], grid[385], grid[386], grid[387], grid[409], grid[411], grid[433], grid[434], grid[435], grid[410]);
evolve8 e411 (grid_evolve[411], grid[386], grid[387], grid[388], grid[410], grid[412], grid[434], grid[435], grid[436], grid[411]);
evolve8 e412 (grid_evolve[412], grid[387], grid[388], grid[389], grid[411], grid[413], grid[435], grid[436], grid[437], grid[412]);
evolve8 e413 (grid_evolve[413], grid[388], grid[389], grid[390], grid[412], grid[414], grid[436], grid[437], grid[438], grid[413]);
evolve8 e414 (grid_evolve[414], grid[389], grid[390], grid[391], grid[413], grid[415], grid[437], grid[438], grid[439], grid[414]);
evolve8 e415 (grid_evolve[415], grid[390], grid[391], grid[392], grid[414], grid[416], grid[438], grid[439], grid[440], grid[415]);
evolve8 e416 (grid_evolve[416], grid[391], grid[392], grid[393], grid[415], grid[417], grid[439], grid[440], grid[441], grid[416]);
evolve8 e417 (grid_evolve[417], grid[392], grid[393], grid[394], grid[416], grid[418], grid[440], grid[441], grid[442], grid[417]);
evolve8 e418 (grid_evolve[418], grid[393], grid[394], grid[395], grid[417], grid[419], grid[441], grid[442], grid[443], grid[418]);
evolve8 e419 (grid_evolve[419], grid[394], grid[395], grid[396], grid[418], grid[420], grid[442], grid[443], grid[444], grid[419]);
evolve8 e420 (grid_evolve[420], grid[395], grid[396], grid[397], grid[419], grid[421], grid[443], grid[444], grid[445], grid[420]);
evolve8 e421 (grid_evolve[421], grid[396], grid[397], grid[398], grid[420], grid[422], grid[444], grid[445], grid[446], grid[421]);
evolve8 e422 (grid_evolve[422], grid[397], grid[398], grid[399], grid[421], grid[423], grid[445], grid[446], grid[447], grid[422]);
evolve8 e423 (grid_evolve[423], grid[398], grid[399], grid[400], grid[422], grid[424], grid[446], grid[447], grid[448], grid[423]);
evolve8 e424 (grid_evolve[424], grid[399], grid[400], grid[401], grid[423], grid[425], grid[447], grid[448], grid[449], grid[424]);
evolve8 e425 (grid_evolve[425], grid[400], grid[401], grid[402], grid[424], grid[426], grid[448], grid[449], grid[450], grid[425]);
evolve8 e426 (grid_evolve[426], grid[401], grid[402], grid[403], grid[425], grid[427], grid[449], grid[450], grid[451], grid[426]);
evolve8 e427 (grid_evolve[427], grid[402], grid[403], grid[404], grid[426], grid[428], grid[450], grid[451], grid[452], grid[427]);
evolve8 e428 (grid_evolve[428], grid[403], grid[404], grid[405], grid[427], grid[429], grid[451], grid[452], grid[453], grid[428]);
evolve8 e429 (grid_evolve[429], grid[404], grid[405], grid[406], grid[428], grid[430], grid[452], grid[453], grid[454], grid[429]);
evolve8 e430 (grid_evolve[430], grid[405], grid[406], grid[407], grid[429], grid[431], grid[453], grid[454], grid[455], grid[430]);
evolve5 e431 (grid_evolve[431], grid[406], grid[407], grid[430], grid[454], grid[455], grid[431]);

evolve5 e432 (grid_evolve[432], grid[408], grid[409], grid[433], grid[456], grid[457], grid[432]);
evolve8 e433 (grid_evolve[433], grid[408], grid[409], grid[410], grid[432], grid[434], grid[456], grid[457], grid[458], grid[433]);
evolve8 e434 (grid_evolve[434], grid[409], grid[410], grid[411], grid[433], grid[435], grid[457], grid[458], grid[459], grid[434]);
evolve8 e435 (grid_evolve[435], grid[410], grid[411], grid[412], grid[434], grid[436], grid[458], grid[459], grid[460], grid[435]);
evolve8 e436 (grid_evolve[436], grid[411], grid[412], grid[413], grid[435], grid[437], grid[459], grid[460], grid[461], grid[436]);
evolve8 e437 (grid_evolve[437], grid[412], grid[413], grid[414], grid[436], grid[438], grid[460], grid[461], grid[462], grid[437]);
evolve8 e438 (grid_evolve[438], grid[413], grid[414], grid[415], grid[437], grid[439], grid[461], grid[462], grid[463], grid[438]);
evolve8 e439 (grid_evolve[439], grid[414], grid[415], grid[416], grid[438], grid[440], grid[462], grid[463], grid[464], grid[439]);
evolve8 e440 (grid_evolve[440], grid[415], grid[416], grid[417], grid[439], grid[441], grid[463], grid[464], grid[465], grid[440]);
evolve8 e441 (grid_evolve[441], grid[416], grid[417], grid[418], grid[440], grid[442], grid[464], grid[465], grid[466], grid[441]);
evolve8 e442 (grid_evolve[442], grid[417], grid[418], grid[419], grid[441], grid[443], grid[465], grid[466], grid[467], grid[442]);
evolve8 e443 (grid_evolve[443], grid[418], grid[419], grid[420], grid[442], grid[444], grid[466], grid[467], grid[468], grid[443]);
evolve8 e444 (grid_evolve[444], grid[419], grid[420], grid[421], grid[443], grid[445], grid[467], grid[468], grid[469], grid[444]);
evolve8 e445 (grid_evolve[445], grid[420], grid[421], grid[422], grid[444], grid[446], grid[468], grid[469], grid[470], grid[445]);
evolve8 e446 (grid_evolve[446], grid[421], grid[422], grid[423], grid[445], grid[447], grid[469], grid[470], grid[471], grid[446]);
evolve8 e447 (grid_evolve[447], grid[422], grid[423], grid[424], grid[446], grid[448], grid[470], grid[471], grid[472], grid[447]);
evolve8 e448 (grid_evolve[448], grid[423], grid[424], grid[425], grid[447], grid[449], grid[471], grid[472], grid[473], grid[448]);
evolve8 e449 (grid_evolve[449], grid[424], grid[425], grid[426], grid[448], grid[450], grid[472], grid[473], grid[474], grid[449]);
evolve8 e450 (grid_evolve[450], grid[425], grid[426], grid[427], grid[449], grid[451], grid[473], grid[474], grid[475], grid[450]);
evolve8 e451 (grid_evolve[451], grid[426], grid[427], grid[428], grid[450], grid[452], grid[474], grid[475], grid[476], grid[451]);
evolve8 e452 (grid_evolve[452], grid[427], grid[428], grid[429], grid[451], grid[453], grid[475], grid[476], grid[477], grid[452]);
evolve8 e453 (grid_evolve[453], grid[428], grid[429], grid[430], grid[452], grid[454], grid[476], grid[477], grid[478], grid[453]);
evolve8 e454 (grid_evolve[454], grid[429], grid[430], grid[431], grid[453], grid[455], grid[477], grid[478], grid[479], grid[454]);
evolve5 e455 (grid_evolve[455], grid[430], grid[431], grid[454], grid[478], grid[479], grid[455]);

evolve5 e456 (grid_evolve[456], grid[432], grid[433], grid[457], grid[480], grid[481], grid[456]);
evolve8 e457 (grid_evolve[457], grid[432], grid[433], grid[434], grid[456], grid[458], grid[480], grid[481], grid[482], grid[457]);
evolve8 e458 (grid_evolve[458], grid[433], grid[434], grid[435], grid[457], grid[459], grid[481], grid[482], grid[483], grid[458]);
evolve8 e459 (grid_evolve[459], grid[434], grid[435], grid[436], grid[458], grid[460], grid[482], grid[483], grid[484], grid[459]);
evolve8 e460 (grid_evolve[460], grid[435], grid[436], grid[437], grid[459], grid[461], grid[483], grid[484], grid[485], grid[460]);
evolve8 e461 (grid_evolve[461], grid[436], grid[437], grid[438], grid[460], grid[462], grid[484], grid[485], grid[486], grid[461]);
evolve8 e462 (grid_evolve[462], grid[437], grid[438], grid[439], grid[461], grid[463], grid[485], grid[486], grid[487], grid[462]);
evolve8 e463 (grid_evolve[463], grid[438], grid[439], grid[440], grid[462], grid[464], grid[486], grid[487], grid[488], grid[463]);
evolve8 e464 (grid_evolve[464], grid[439], grid[440], grid[441], grid[463], grid[465], grid[487], grid[488], grid[489], grid[464]);
evolve8 e465 (grid_evolve[465], grid[440], grid[441], grid[442], grid[464], grid[466], grid[488], grid[489], grid[490], grid[465]);
evolve8 e466 (grid_evolve[466], grid[441], grid[442], grid[443], grid[465], grid[467], grid[489], grid[490], grid[491], grid[466]);
evolve8 e467 (grid_evolve[467], grid[442], grid[443], grid[444], grid[466], grid[468], grid[490], grid[491], grid[492], grid[467]);
evolve8 e468 (grid_evolve[468], grid[443], grid[444], grid[445], grid[467], grid[469], grid[491], grid[492], grid[493], grid[468]);
evolve8 e469 (grid_evolve[469], grid[444], grid[445], grid[446], grid[468], grid[470], grid[492], grid[493], grid[494], grid[469]);
evolve8 e470 (grid_evolve[470], grid[445], grid[446], grid[447], grid[469], grid[471], grid[493], grid[494], grid[495], grid[470]);
evolve8 e471 (grid_evolve[471], grid[446], grid[447], grid[448], grid[470], grid[472], grid[494], grid[495], grid[496], grid[471]);
evolve8 e472 (grid_evolve[472], grid[447], grid[448], grid[449], grid[471], grid[473], grid[495], grid[496], grid[497], grid[472]);
evolve8 e473 (grid_evolve[473], grid[448], grid[449], grid[450], grid[472], grid[474], grid[496], grid[497], grid[498], grid[473]);
evolve8 e474 (grid_evolve[474], grid[449], grid[450], grid[451], grid[473], grid[475], grid[497], grid[498], grid[499], grid[474]);
evolve8 e475 (grid_evolve[475], grid[450], grid[451], grid[452], grid[474], grid[476], grid[498], grid[499], grid[500], grid[475]);
evolve8 e476 (grid_evolve[476], grid[451], grid[452], grid[453], grid[475], grid[477], grid[499], grid[500], grid[501], grid[476]);
evolve8 e477 (grid_evolve[477], grid[452], grid[453], grid[454], grid[476], grid[478], grid[500], grid[501], grid[502], grid[477]);
evolve8 e478 (grid_evolve[478], grid[453], grid[454], grid[455], grid[477], grid[479], grid[501], grid[502], grid[503], grid[478]);
evolve5 e479 (grid_evolve[479], grid[454], grid[455], grid[478], grid[502], grid[503], grid[479]);

evolve5 e480 (grid_evolve[480], grid[456], grid[457], grid[481], grid[504], grid[505], grid[480]);
evolve8 e481 (grid_evolve[481], grid[456], grid[457], grid[458], grid[480], grid[482], grid[504], grid[505], grid[506], grid[481]);
evolve8 e482 (grid_evolve[482], grid[457], grid[458], grid[459], grid[481], grid[483], grid[505], grid[506], grid[507], grid[482]);
evolve8 e483 (grid_evolve[483], grid[458], grid[459], grid[460], grid[482], grid[484], grid[506], grid[507], grid[508], grid[483]);
evolve8 e484 (grid_evolve[484], grid[459], grid[460], grid[461], grid[483], grid[485], grid[507], grid[508], grid[509], grid[484]);
evolve8 e485 (grid_evolve[485], grid[460], grid[461], grid[462], grid[484], grid[486], grid[508], grid[509], grid[510], grid[485]);
evolve8 e486 (grid_evolve[486], grid[461], grid[462], grid[463], grid[485], grid[487], grid[509], grid[510], grid[511], grid[486]);
evolve8 e487 (grid_evolve[487], grid[462], grid[463], grid[464], grid[486], grid[488], grid[510], grid[511], grid[512], grid[487]);
evolve8 e488 (grid_evolve[488], grid[463], grid[464], grid[465], grid[487], grid[489], grid[511], grid[512], grid[513], grid[488]);
evolve8 e489 (grid_evolve[489], grid[464], grid[465], grid[466], grid[488], grid[490], grid[512], grid[513], grid[514], grid[489]);
evolve8 e490 (grid_evolve[490], grid[465], grid[466], grid[467], grid[489], grid[491], grid[513], grid[514], grid[515], grid[490]);
evolve8 e491 (grid_evolve[491], grid[466], grid[467], grid[468], grid[490], grid[492], grid[514], grid[515], grid[516], grid[491]);
evolve8 e492 (grid_evolve[492], grid[467], grid[468], grid[469], grid[491], grid[493], grid[515], grid[516], grid[517], grid[492]);
evolve8 e493 (grid_evolve[493], grid[468], grid[469], grid[470], grid[492], grid[494], grid[516], grid[517], grid[518], grid[493]);
evolve8 e494 (grid_evolve[494], grid[469], grid[470], grid[471], grid[493], grid[495], grid[517], grid[518], grid[519], grid[494]);
evolve8 e495 (grid_evolve[495], grid[470], grid[471], grid[472], grid[494], grid[496], grid[518], grid[519], grid[520], grid[495]);
evolve8 e496 (grid_evolve[496], grid[471], grid[472], grid[473], grid[495], grid[497], grid[519], grid[520], grid[521], grid[496]);
evolve8 e497 (grid_evolve[497], grid[472], grid[473], grid[474], grid[496], grid[498], grid[520], grid[521], grid[522], grid[497]);
evolve8 e498 (grid_evolve[498], grid[473], grid[474], grid[475], grid[497], grid[499], grid[521], grid[522], grid[523], grid[498]);
evolve8 e499 (grid_evolve[499], grid[474], grid[475], grid[476], grid[498], grid[500], grid[522], grid[523], grid[524], grid[499]);
evolve8 e500 (grid_evolve[500], grid[475], grid[476], grid[477], grid[499], grid[501], grid[523], grid[524], grid[525], grid[500]);
evolve8 e501 (grid_evolve[501], grid[476], grid[477], grid[478], grid[500], grid[502], grid[524], grid[525], grid[526], grid[501]);
evolve8 e502 (grid_evolve[502], grid[477], grid[478], grid[479], grid[501], grid[503], grid[525], grid[526], grid[527], grid[502]);
evolve5 e503 (grid_evolve[503], grid[478], grid[479], grid[502], grid[526], grid[527], grid[503]);

evolve5 e504 (grid_evolve[504], grid[480], grid[481], grid[505], grid[528], grid[529], grid[504]);
evolve8 e505 (grid_evolve[505], grid[480], grid[481], grid[482], grid[504], grid[506], grid[528], grid[529], grid[530], grid[505]);
evolve8 e506 (grid_evolve[506], grid[481], grid[482], grid[483], grid[505], grid[507], grid[529], grid[530], grid[531], grid[506]);
evolve8 e507 (grid_evolve[507], grid[482], grid[483], grid[484], grid[506], grid[508], grid[530], grid[531], grid[532], grid[507]);
evolve8 e508 (grid_evolve[508], grid[483], grid[484], grid[485], grid[507], grid[509], grid[531], grid[532], grid[533], grid[508]);
evolve8 e509 (grid_evolve[509], grid[484], grid[485], grid[486], grid[508], grid[510], grid[532], grid[533], grid[534], grid[509]);
evolve8 e510 (grid_evolve[510], grid[485], grid[486], grid[487], grid[509], grid[511], grid[533], grid[534], grid[535], grid[510]);
evolve8 e511 (grid_evolve[511], grid[486], grid[487], grid[488], grid[510], grid[512], grid[534], grid[535], grid[536], grid[511]);
evolve8 e512 (grid_evolve[512], grid[487], grid[488], grid[489], grid[511], grid[513], grid[535], grid[536], grid[537], grid[512]);
evolve8 e513 (grid_evolve[513], grid[488], grid[489], grid[490], grid[512], grid[514], grid[536], grid[537], grid[538], grid[513]);
evolve8 e514 (grid_evolve[514], grid[489], grid[490], grid[491], grid[513], grid[515], grid[537], grid[538], grid[539], grid[514]);
evolve8 e515 (grid_evolve[515], grid[490], grid[491], grid[492], grid[514], grid[516], grid[538], grid[539], grid[540], grid[515]);
evolve8 e516 (grid_evolve[516], grid[491], grid[492], grid[493], grid[515], grid[517], grid[539], grid[540], grid[541], grid[516]);
evolve8 e517 (grid_evolve[517], grid[492], grid[493], grid[494], grid[516], grid[518], grid[540], grid[541], grid[542], grid[517]);
evolve8 e518 (grid_evolve[518], grid[493], grid[494], grid[495], grid[517], grid[519], grid[541], grid[542], grid[543], grid[518]);
evolve8 e519 (grid_evolve[519], grid[494], grid[495], grid[496], grid[518], grid[520], grid[542], grid[543], grid[544], grid[519]);
evolve8 e520 (grid_evolve[520], grid[495], grid[496], grid[497], grid[519], grid[521], grid[543], grid[544], grid[545], grid[520]);
evolve8 e521 (grid_evolve[521], grid[496], grid[497], grid[498], grid[520], grid[522], grid[544], grid[545], grid[546], grid[521]);
evolve8 e522 (grid_evolve[522], grid[497], grid[498], grid[499], grid[521], grid[523], grid[545], grid[546], grid[547], grid[522]);
evolve8 e523 (grid_evolve[523], grid[498], grid[499], grid[500], grid[522], grid[524], grid[546], grid[547], grid[548], grid[523]);
evolve8 e524 (grid_evolve[524], grid[499], grid[500], grid[501], grid[523], grid[525], grid[547], grid[548], grid[549], grid[524]);
evolve8 e525 (grid_evolve[525], grid[500], grid[501], grid[502], grid[524], grid[526], grid[548], grid[549], grid[550], grid[525]);
evolve8 e526 (grid_evolve[526], grid[501], grid[502], grid[503], grid[525], grid[527], grid[549], grid[550], grid[551], grid[526]);
evolve5 e527 (grid_evolve[527], grid[502], grid[503], grid[526], grid[550], grid[551], grid[527]);

evolve5 e528 (grid_evolve[528], grid[504], grid[505], grid[529], grid[552], grid[553], grid[528]);
evolve8 e529 (grid_evolve[529], grid[504], grid[505], grid[506], grid[528], grid[530], grid[552], grid[553], grid[554], grid[529]);
evolve8 e530 (grid_evolve[530], grid[505], grid[506], grid[507], grid[529], grid[531], grid[553], grid[554], grid[555], grid[530]);
evolve8 e531 (grid_evolve[531], grid[506], grid[507], grid[508], grid[530], grid[532], grid[554], grid[555], grid[556], grid[531]);
evolve8 e532 (grid_evolve[532], grid[507], grid[508], grid[509], grid[531], grid[533], grid[555], grid[556], grid[557], grid[532]);
evolve8 e533 (grid_evolve[533], grid[508], grid[509], grid[510], grid[532], grid[534], grid[556], grid[557], grid[558], grid[533]);
evolve8 e534 (grid_evolve[534], grid[509], grid[510], grid[511], grid[533], grid[535], grid[557], grid[558], grid[559], grid[534]);
evolve8 e535 (grid_evolve[535], grid[510], grid[511], grid[512], grid[534], grid[536], grid[558], grid[559], grid[560], grid[535]);
evolve8 e536 (grid_evolve[536], grid[511], grid[512], grid[513], grid[535], grid[537], grid[559], grid[560], grid[561], grid[536]);
evolve8 e537 (grid_evolve[537], grid[512], grid[513], grid[514], grid[536], grid[538], grid[560], grid[561], grid[562], grid[537]);
evolve8 e538 (grid_evolve[538], grid[513], grid[514], grid[515], grid[537], grid[539], grid[561], grid[562], grid[563], grid[538]);
evolve8 e539 (grid_evolve[539], grid[514], grid[515], grid[516], grid[538], grid[540], grid[562], grid[563], grid[564], grid[539]);
evolve8 e540 (grid_evolve[540], grid[515], grid[516], grid[517], grid[539], grid[541], grid[563], grid[564], grid[565], grid[540]);
evolve8 e541 (grid_evolve[541], grid[516], grid[517], grid[518], grid[540], grid[542], grid[564], grid[565], grid[566], grid[541]);
evolve8 e542 (grid_evolve[542], grid[517], grid[518], grid[519], grid[541], grid[543], grid[565], grid[566], grid[567], grid[542]);
evolve8 e543 (grid_evolve[543], grid[518], grid[519], grid[520], grid[542], grid[544], grid[566], grid[567], grid[568], grid[543]);
evolve8 e544 (grid_evolve[544], grid[519], grid[520], grid[521], grid[543], grid[545], grid[567], grid[568], grid[569], grid[544]);
evolve8 e545 (grid_evolve[545], grid[520], grid[521], grid[522], grid[544], grid[546], grid[568], grid[569], grid[570], grid[545]);
evolve8 e546 (grid_evolve[546], grid[521], grid[522], grid[523], grid[545], grid[547], grid[569], grid[570], grid[571], grid[546]);
evolve8 e547 (grid_evolve[547], grid[522], grid[523], grid[524], grid[546], grid[548], grid[570], grid[571], grid[572], grid[547]);
evolve8 e548 (grid_evolve[548], grid[523], grid[524], grid[525], grid[547], grid[549], grid[571], grid[572], grid[573], grid[548]);
evolve8 e549 (grid_evolve[549], grid[524], grid[525], grid[526], grid[548], grid[550], grid[572], grid[573], grid[574], grid[549]);
evolve8 e550 (grid_evolve[550], grid[525], grid[526], grid[527], grid[549], grid[551], grid[573], grid[574], grid[575], grid[550]);
evolve5 e551 (grid_evolve[551], grid[526], grid[527], grid[550], grid[574], grid[575], grid[551]);

evolve3 e552 (grid_evolve[552], grid[528], grid[529], grid[553], grid[552]);
evolve5 e553 (grid_evolve[553], grid[528], grid[529], grid[530], grid[552], grid[554], grid[553]);
evolve5 e554 (grid_evolve[554], grid[529], grid[530], grid[531], grid[553], grid[555], grid[554]);
evolve5 e555 (grid_evolve[555], grid[530], grid[531], grid[532], grid[554], grid[556], grid[555]);
evolve5 e556 (grid_evolve[556], grid[531], grid[532], grid[533], grid[555], grid[557], grid[556]);
evolve5 e557 (grid_evolve[557], grid[532], grid[533], grid[534], grid[556], grid[558], grid[557]);
evolve5 e558 (grid_evolve[558], grid[533], grid[534], grid[535], grid[557], grid[559], grid[558]);
evolve5 e559 (grid_evolve[559], grid[534], grid[535], grid[536], grid[558], grid[560], grid[559]);
evolve5 e560 (grid_evolve[560], grid[535], grid[536], grid[537], grid[559], grid[561], grid[560]);
evolve5 e561 (grid_evolve[561], grid[536], grid[537], grid[538], grid[560], grid[562], grid[561]);
evolve5 e562 (grid_evolve[562], grid[537], grid[538], grid[539], grid[561], grid[563], grid[562]);
evolve5 e563 (grid_evolve[563], grid[538], grid[539], grid[540], grid[562], grid[564], grid[563]);
evolve5 e564 (grid_evolve[564], grid[539], grid[540], grid[541], grid[563], grid[565], grid[564]);
evolve5 e565 (grid_evolve[565], grid[540], grid[541], grid[542], grid[564], grid[566], grid[565]);
evolve5 e566 (grid_evolve[566], grid[541], grid[542], grid[543], grid[565], grid[567], grid[566]);
evolve5 e567 (grid_evolve[567], grid[542], grid[543], grid[544], grid[566], grid[568], grid[567]);
evolve5 e568 (grid_evolve[568], grid[543], grid[544], grid[545], grid[567], grid[569], grid[568]);
evolve5 e569 (grid_evolve[569], grid[544], grid[545], grid[546], grid[568], grid[570], grid[569]);
evolve5 e570 (grid_evolve[570], grid[545], grid[546], grid[547], grid[569], grid[571], grid[570]);
evolve5 e571 (grid_evolve[571], grid[546], grid[547], grid[548], grid[570], grid[572], grid[571]);
evolve5 e572 (grid_evolve[572], grid[547], grid[548], grid[549], grid[571], grid[573], grid[572]);
evolve5 e573 (grid_evolve[573], grid[548], grid[549], grid[550], grid[572], grid[574], grid[573]);
evolve5 e574 (grid_evolve[574], grid[549], grid[550], grid[551], grid[573], grid[575], grid[574]);
evolve3 e575 (grid_evolve[575], grid[550], grid[551], grid[574], grid[575]);
 
endmodule // top


module evolve3 (next_state, vector1, vector2, vector3, current_state);
	
   input logic  vector1;
   input logic  vector2;
   input logic  vector3;
   input logic  current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve3

module evolve5 (next_state, vector1, vector2, vector3, 
		vector4, vector5, current_state);
   
   input logic     vector1;
   input logic 	 vector2;
   input logic 	 vector3;
   input logic 	 vector4;
   input logic 	 vector5;
   input logic 	 current_state;
   output logic    next_state;
   
   logic [3:0] 	 sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + vector5;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve5


module evolve8 (next_state, vector1, vector2, vector3, 
		vector4, vector5, vector6, 
		vector7, vector8, current_state);
   
   input logic 	vector1;
   input logic 	vector2;
   input logic 	vector3;
   input logic 	vector4;
   input logic 	vector5;
	
   input logic 	vector6;
   input logic 	vector7;
   input logic 	vector8;
   input logic 	current_state;
   output logic   next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + 
		vector5 + vector6 + vector7 + vector8;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve8


module rules (pop_count, current_state, next_state);
   
   input logic [3:0] pop_count;
   input logic 	     current_state;
   output logic      next_state;
   
   assign next_state = (pop_count == 2 & current_state) | pop_count == 3;
   
endmodule // rules